library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Seed is
	
	constant 

end package ; -- Seed 