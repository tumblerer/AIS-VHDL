LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.test_core;
USE work.project_pak.ALL;
USE work.utility.ALL;

USE std.textio.ALL;
use ieee.std_logic_textio.all;
use work.Pack.all;


ENTITY test_core_test_bench IS

END ENTITY test_core_test_bench;

ARCHITECTURE test_bench OF test_core_test_bench IS

SIGNAL SYS_CLK, SYS_RST : std_logic := '0';

signal INPUT_1 : std_logic_vector(31 downto 0) := "00000000000000000000000000000110";
signal INPUT_2 : std_logic_vector(31 downto 0) := "00000000000000000000000000010100";
signal INPUT_3 : std_logic_vector(31 downto 0) := "00111111111100000000000000000000";
signal INPUT_4 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_5 : std_logic_vector(31 downto 0) := "00111111101110011001100110011001";
signal INPUT_6 : std_logic_vector(31 downto 0) := "10011001100110011001100110011010";
signal INPUT_7 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_8 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_9 : std_logic_vector(31 downto 0) := "00111111111100000000000000000000";
signal INPUT_10 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_11 : std_logic_vector(31 downto 0) := "00111111101010011001100110011001";
signal INPUT_12 : std_logic_vector(31 downto 0) := "10011001100110011001100110011010";
signal INPUT_13 : std_logic_vector(31 downto 0) := "00111111110001010101010101010101";
signal INPUT_14 : std_logic_vector(31 downto 0) := "01010101010101010101010101010101";
signal INPUT_15 : std_logic_vector(31 downto 0) := "00111111110101010101010101010101";
signal INPUT_16 : std_logic_vector(31 downto 0) := "01010101010101010101010101010101";
signal INPUT_17 : std_logic_vector(31 downto 0) := "00111111111000000000000000000000";
signal INPUT_18 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_19 : std_logic_vector(31 downto 0) := "00111111111001010101010101010101";
signal INPUT_20 : std_logic_vector(31 downto 0) := "01010101010101010101010101010101";
signal INPUT_21 : std_logic_vector(31 downto 0) := "00111111111010101010101010101010";
signal INPUT_22 : std_logic_vector(31 downto 0) := "10101010101010101010101010101011";
signal INPUT_23 : std_logic_vector(31 downto 0) := "00111111111100000000000000000000";
signal INPUT_24 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_25 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_26 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_27 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_28 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_29 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_30 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_31 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_32 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_33 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_34 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_35 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_36 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_37 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_38 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_39 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_40 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_41 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_42 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_43 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_44 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_45 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_46 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_47 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_48 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_49 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_50 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_51 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_52 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_53 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_54 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_55 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_56 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_57 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_58 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_59 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_60 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_61 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_62 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_63 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_64 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_65 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_66 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_67 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_68 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_69 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_70 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_71 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_72 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_73 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_74 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_75 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_76 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_77 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_78 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_79 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_80 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_81 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_82 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_83 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_84 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_85 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_86 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_87 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_88 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_89 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_90 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_91 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_92 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_93 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_94 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_95 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_96 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_97 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_98 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_99 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_100 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_101 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_102 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_103 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_104 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_105 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_106 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_107 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_108 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_109 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_110 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_111 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_112 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_113 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_114 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_115 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_116 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_117 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_118 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_119 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_120 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_121 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_122 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_123 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_124 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_125 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_126 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_127 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_128 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_129 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_130 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_131 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_132 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_133 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_134 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_135 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_136 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_137 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_138 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_139 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_140 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_141 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_142 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_143 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_144 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_145 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_146 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_147 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_148 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_149 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_150 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_151 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_152 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_153 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_154 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_155 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_156 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_157 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_158 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_159 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_160 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_161 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_162 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_163 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_164 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_165 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_166 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_167 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_168 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_169 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_170 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_171 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_172 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_173 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_174 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_175 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_176 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_177 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_178 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_179 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_180 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_181 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_182 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_183 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_184 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_185 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_186 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_187 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_188 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_189 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_190 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_191 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_192 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_193 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_194 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_195 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_196 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_197 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_198 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_199 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_200 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_201 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_202 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_203 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_204 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_205 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_206 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_207 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_208 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_209 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_210 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_211 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_212 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_213 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_214 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_215 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_216 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_217 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_218 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_219 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_220 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_221 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_222 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_223 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_224 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_225 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_226 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_227 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_228 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_229 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_230 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_231 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_232 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_233 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_234 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_235 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_236 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_237 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_238 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_239 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_240 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_241 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_242 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_243 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_244 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_245 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_246 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_247 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_248 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_249 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_250 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_251 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_252 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_253 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_254 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_255 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_256 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_257 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_258 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_259 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_260 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_261 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_262 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_263 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_264 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_265 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_266 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_267 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_268 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_269 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_270 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_271 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_272 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_273 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_274 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_275 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_276 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_277 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_278 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_279 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_280 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_281 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_282 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_283 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_284 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_285 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_286 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_287 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_288 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_289 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_290 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_291 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_292 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_293 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_294 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_295 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_296 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_297 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_298 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_299 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_300 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_301 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_302 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_303 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_304 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_305 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_306 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_307 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_308 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_309 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_310 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_311 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_312 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_313 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_314 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_315 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_316 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_317 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_318 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_319 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_320 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_321 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_322 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_323 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_324 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_325 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_326 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_327 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_328 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_329 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_330 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_331 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_332 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_333 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_334 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_335 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_336 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_337 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_338 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_339 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_340 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_341 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_342 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_343 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_344 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_345 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_346 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_347 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_348 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_349 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_350 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_351 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_352 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_353 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_354 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_355 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_356 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_357 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_358 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_359 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_360 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_361 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_362 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_363 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_364 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_365 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_366 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_367 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_368 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_369 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_370 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_371 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_372 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_373 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_374 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_375 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_376 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_377 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_378 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_379 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_380 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_381 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_382 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_383 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_384 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_385 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_386 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_387 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_388 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_389 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_390 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_391 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_392 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_393 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_394 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_395 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_396 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_397 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_398 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_399 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_400 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_401 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_402 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_403 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_404 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_405 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_406 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_407 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_408 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_409 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_410 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_411 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_412 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_413 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_414 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_415 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_416 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_417 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_418 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_419 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_420 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_421 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_422 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_423 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_424 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_425 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_426 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_427 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_428 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_429 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_430 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_431 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_432 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_433 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_434 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_435 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_436 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_437 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_438 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_439 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_440 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_441 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_442 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_443 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_444 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_445 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_446 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_447 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_448 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_449 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_450 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_451 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_452 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_453 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_454 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_455 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_456 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_457 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_458 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_459 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_460 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_461 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_462 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_463 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_464 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_465 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_466 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_467 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_468 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_469 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_470 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_471 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_472 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_473 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_474 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_475 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_476 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_477 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_478 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_479 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_480 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_481 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_482 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_483 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_484 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_485 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_486 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_487 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_488 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_489 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_490 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_491 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_492 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_493 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_494 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_495 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_496 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_497 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_498 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_499 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_500 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_501 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_502 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_503 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_504 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_505 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_506 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_507 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_508 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_509 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_510 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_511 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_512 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_513 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_514 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_515 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_516 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_517 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_518 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_519 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_520 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_521 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_522 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_523 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_524 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_525 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_526 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_527 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_528 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_529 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_530 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_531 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_532 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_533 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_534 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_535 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_536 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_537 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_538 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_539 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_540 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_541 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_542 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_543 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_544 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_545 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_546 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_547 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_548 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_549 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_550 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_551 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_552 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_553 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_554 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_555 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_556 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_557 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_558 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_559 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_560 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_561 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_562 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_563 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_564 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_565 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_566 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_567 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_568 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_569 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_570 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_571 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_572 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_573 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_574 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_575 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_576 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_577 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_578 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_579 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_580 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_581 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_582 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_583 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_584 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_585 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_586 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_587 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_588 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_589 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_590 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_591 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_592 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_593 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_594 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_595 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_596 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_597 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_598 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_599 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_600 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_601 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_602 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_603 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_604 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_605 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_606 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_607 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_608 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_609 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_610 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_611 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_612 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_613 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_614 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
signal INPUT_615 : std_logic_vector(31 downto 0) := "00111111111010100001001000110111";
signal INPUT_616 : std_logic_vector(31 downto 0) := "01101000100010101011101001111011";
signal INPUT_617 : std_logic_vector(31 downto 0) := "00111111111011001111110000111111";
signal INPUT_618 : std_logic_vector(31 downto 0) := "01011111010101110000110001111101";
signal INPUT_619 : std_logic_vector(31 downto 0) := "00111111110000000100000100011010";
signal INPUT_620 : std_logic_vector(31 downto 0) := "10011111100000000111101101111100";
signal INPUT_621 : std_logic_vector(31 downto 0) := "00111111111011010011101001100000";
signal INPUT_622 : std_logic_vector(31 downto 0) := "00000000111000100101011010111111";
signal INPUT_623 : std_logic_vector(31 downto 0) := "00111111111001000011110001001001";
signal INPUT_624 : std_logic_vector(31 downto 0) := "01110101001110111001000000100100";
signal INPUT_625 : std_logic_vector(31 downto 0) := "00111111101110001111100001101000";
signal INPUT_626 : std_logic_vector(31 downto 0) := "01110001100000101101010011000000";
signal INPUT_627 : std_logic_vector(31 downto 0) := "00111111110100011101001011101010";
signal INPUT_628 : std_logic_vector(31 downto 0) := "00110001100000011100111001101000";
signal INPUT_629 : std_logic_vector(31 downto 0) := "00111111111000011000000000001101";
signal INPUT_630 : std_logic_vector(31 downto 0) := "10101011111110001011010111100000";
signal INPUT_631 : std_logic_vector(31 downto 0) := "00111111111011101010001111100101";
signal INPUT_632 : std_logic_vector(31 downto 0) := "01011111111111000110000001011011";
signal INPUT_633 : std_logic_vector(31 downto 0) := "00111111111011101110000001011101";
signal INPUT_634 : std_logic_vector(31 downto 0) := "11101011110111101110101101101011";
signal INPUT_635 : std_logic_vector(31 downto 0) := "00111111110001000010110010101010";
signal INPUT_636 : std_logic_vector(31 downto 0) := "01011011100111010000100101010000";
signal INPUT_637 : std_logic_vector(31 downto 0) := "00111111111011110000111100011000";
signal INPUT_638 : std_logic_vector(31 downto 0) := "10010111111011001010100000000100";
signal INPUT_639 : std_logic_vector(31 downto 0) := "00111111111011101010000100011100";
signal INPUT_640 : std_logic_vector(31 downto 0) := "10010100011100000111111110011001";
signal INPUT_641 : std_logic_vector(31 downto 0) := "00111111110111110001000001100101";
signal INPUT_642 : std_logic_vector(31 downto 0) := "00000110011000101000010101010010";
signal INPUT_643 : std_logic_vector(31 downto 0) := "00111111111010011001101111100101";
signal INPUT_644 : std_logic_vector(31 downto 0) := "11001001001100000010100001111100";
signal INPUT_645 : std_logic_vector(31 downto 0) := "00111111110000100010100101010100";
signal INPUT_646 : std_logic_vector(31 downto 0) := "11100000000100111001011111011000";
signal INPUT_647 : std_logic_vector(31 downto 0) := "00111111110110101111111000100011";
signal INPUT_648 : std_logic_vector(31 downto 0) := "00001000111001100101001111001010";
signal INPUT_649 : std_logic_vector(31 downto 0) := "00111111111011010100110110110100";
signal INPUT_650 : std_logic_vector(31 downto 0) := "10010110100011110001111000100000";
signal INPUT_651 : std_logic_vector(31 downto 0) := "00111111111010010101100111000011";
signal INPUT_652 : std_logic_vector(31 downto 0) := "00101111100000111000001101010010";
signal INPUT_653 : std_logic_vector(31 downto 0) := "00111111111011101011010000101001";
signal INPUT_654 : std_logic_vector(31 downto 0) := "01110110000000111100000000100110";



SIGNAL OUTPUT : std_logic_vector(32 - 1 DOWNTO 0);
SIGNAL OUTPUT_2 : std_logic_vector(32 - 1 DOWNTO 0);

SIGNAL VALID : std_logic := '0';

SIGNAL START : std_logic := '0';

SIGNAL RUNTIME : std_logic_vector(32 - 1 DOWNTO 0);

SIGNAL FINISHED : std_logic := '0';

SIGNAL BUSY : std_logic := '0';

SIGNAL OUTPUT_CYCLE : std_logic_vector(32 - 1  DOWNTO 0);

SIGNAL i : integer := 0;

signal steps, runs : std_logic_vector(31 downto 0);

BEGIN

DUT : ENTITY work.test_core
  GENERIC MAP(
    C_SIMPBUS_AWIDTH  => 32
  )
  PORT MAP(
    SYS_CLK     => SYS_CLK,
    SYS_RST     => SYS_RST,
    INPUT_1       => INPUT_1,
    INPUT_2       => INPUT_2,
    INPUT_3       => INPUT_3,
    INPUT_4       => INPUT_4,
    INPUT_5       => INPUT_5,
    INPUT_6       => INPUT_6,
    INPUT_7       => INPUT_7,
    INPUT_8       => INPUT_8,
    INPUT_9       => INPUT_9,
    INPUT_10      => INPUT_10,
    INPUT_11      => INPUT_11,
    INPUT_12      => INPUT_12,
    INPUT_13      => INPUT_13,
    INPUT_14      => INPUT_14,
    INPUT_15      => INPUT_15,
    INPUT_16      => INPUT_16,
    INPUT_17      => INPUT_17,
    INPUT_18      => INPUT_18,
    INPUT_19      => INPUT_19,
    INPUT_20      => INPUT_20,
    INPUT_21      => INPUT_21,
    INPUT_22      => INPUT_22,
    INPUT_23      => INPUT_23,
    INPUT_24      => INPUT_24,
    INPUT_25      => INPUT_25,
    INPUT_26      => INPUT_26,
    INPUT_27      => INPUT_27,
    INPUT_28      => INPUT_28,
    INPUT_29      => INPUT_29,
    INPUT_30      => INPUT_30,
    INPUT_31      => INPUT_31,
    INPUT_32      => INPUT_32,
    INPUT_33      => INPUT_33,
    INPUT_34      => INPUT_34,
    INPUT_35      => INPUT_35,
    INPUT_36      => INPUT_36,
    INPUT_37      => INPUT_37,
    INPUT_38      => INPUT_38,
    INPUT_39      => INPUT_39,
    INPUT_40      => INPUT_40,
    INPUT_41      => INPUT_41,
    INPUT_42      => INPUT_42,
    INPUT_43      => INPUT_43,
    INPUT_44      => INPUT_44,
    INPUT_45      => INPUT_45,
    INPUT_46      => INPUT_46,
    INPUT_47      => INPUT_47,
    INPUT_48      => INPUT_48,
    INPUT_49      => INPUT_49,
    INPUT_50      => INPUT_50,
    INPUT_51      => INPUT_51,
    INPUT_52      => INPUT_52,
    INPUT_53      => INPUT_53,
    INPUT_54      => INPUT_54,
    INPUT_55      => INPUT_55,
    INPUT_56      => INPUT_56,
    INPUT_57      => INPUT_57,
    INPUT_58      => INPUT_58,
    INPUT_59      => INPUT_59,
    INPUT_60      => INPUT_60,
    INPUT_61      => INPUT_61,
    INPUT_62      => INPUT_62,
    INPUT_63      => INPUT_63,
    INPUT_64      => INPUT_64,
    INPUT_65      => INPUT_65,
    INPUT_66      => INPUT_66,
    INPUT_67      => INPUT_67,
    INPUT_68      => INPUT_68,
    INPUT_69      => INPUT_69,
    INPUT_70      => INPUT_70,
    INPUT_71      => INPUT_71,
    INPUT_72      => INPUT_72,
    INPUT_73      => INPUT_73,
    INPUT_74      => INPUT_74,
    INPUT_75      => INPUT_75,
    INPUT_76      => INPUT_76,
    INPUT_77      => INPUT_77,
    INPUT_78      => INPUT_78,
    INPUT_79      => INPUT_79,
    INPUT_80      => INPUT_80,
    INPUT_81      => INPUT_81,
    INPUT_82      => INPUT_82,
    INPUT_83      => INPUT_83,
    INPUT_84      => INPUT_84,
    INPUT_85      => INPUT_85,
    INPUT_86      => INPUT_86,
    INPUT_87      => INPUT_87,
    INPUT_88      => INPUT_88,
    INPUT_89      => INPUT_89,
    INPUT_90      => INPUT_90,
    INPUT_91      => INPUT_91,
    INPUT_92      => INPUT_92,
    INPUT_93      => INPUT_93,
    INPUT_94      => INPUT_94,
    INPUT_95      => INPUT_95,
    INPUT_96      => INPUT_96,
    INPUT_97      => INPUT_97,
    INPUT_98      => INPUT_98,
    INPUT_99      => INPUT_99,
    INPUT_100       => INPUT_100,
    INPUT_101       => INPUT_101,
    INPUT_102       => INPUT_102,
    INPUT_103       => INPUT_103,
    INPUT_104       => INPUT_104,
    INPUT_105       => INPUT_105,
    INPUT_106       => INPUT_106,
    INPUT_107       => INPUT_107,
    INPUT_108       => INPUT_108,
    INPUT_109       => INPUT_109,
    INPUT_110       => INPUT_110,
    INPUT_111       => INPUT_111,
    INPUT_112       => INPUT_112,
    INPUT_113       => INPUT_113,
    INPUT_114       => INPUT_114,
    INPUT_115       => INPUT_115,
    INPUT_116       => INPUT_116,
    INPUT_117       => INPUT_117,
    INPUT_118       => INPUT_118,
    INPUT_119       => INPUT_119,
    INPUT_120       => INPUT_120,
    INPUT_121       => INPUT_121,
    INPUT_122       => INPUT_122,
    INPUT_123       => INPUT_123,
    INPUT_124       => INPUT_124,
    INPUT_125       => INPUT_125,
    INPUT_126       => INPUT_126,
    INPUT_127       => INPUT_127,
    INPUT_128       => INPUT_128,
    INPUT_129       => INPUT_129,
    INPUT_130       => INPUT_130,
    INPUT_131       => INPUT_131,
    INPUT_132       => INPUT_132,
    INPUT_133       => INPUT_133,
    INPUT_134       => INPUT_134,
    INPUT_135       => INPUT_135,
    INPUT_136       => INPUT_136,
    INPUT_137       => INPUT_137,
    INPUT_138       => INPUT_138,
    INPUT_139       => INPUT_139,
    INPUT_140       => INPUT_140,
    INPUT_141       => INPUT_141,
    INPUT_142       => INPUT_142,
    INPUT_143       => INPUT_143,
    INPUT_144       => INPUT_144,
    INPUT_145       => INPUT_145,
    INPUT_146       => INPUT_146,
    INPUT_147       => INPUT_147,
    INPUT_148       => INPUT_148,
    INPUT_149       => INPUT_149,
    INPUT_150       => INPUT_150,
    INPUT_151       => INPUT_151,
    INPUT_152       => INPUT_152,
    INPUT_153       => INPUT_153,
    INPUT_154       => INPUT_154,
    INPUT_155       => INPUT_155,
    INPUT_156       => INPUT_156,
    INPUT_157       => INPUT_157,
    INPUT_158       => INPUT_158,
    INPUT_159       => INPUT_159,
    INPUT_160       => INPUT_160,
    INPUT_161       => INPUT_161,
    INPUT_162       => INPUT_162,
    INPUT_163       => INPUT_163,
    INPUT_164       => INPUT_164,
    INPUT_165       => INPUT_165,
    INPUT_166       => INPUT_166,
    INPUT_167       => INPUT_167,
    INPUT_168       => INPUT_168,
    INPUT_169       => INPUT_169,
    INPUT_170       => INPUT_170,
    INPUT_171       => INPUT_171,
    INPUT_172       => INPUT_172,
    INPUT_173       => INPUT_173,
    INPUT_174       => INPUT_174,
    INPUT_175       => INPUT_175,
    INPUT_176       => INPUT_176,
    INPUT_177       => INPUT_177,
    INPUT_178       => INPUT_178,
    INPUT_179       => INPUT_179,
    INPUT_180       => INPUT_180,
    INPUT_181       => INPUT_181,
    INPUT_182       => INPUT_182,
    INPUT_183       => INPUT_183,
    INPUT_184       => INPUT_184,
    INPUT_185       => INPUT_185,
    INPUT_186       => INPUT_186,
    INPUT_187       => INPUT_187,
    INPUT_188       => INPUT_188,
    INPUT_189       => INPUT_189,
    INPUT_190       => INPUT_190,
    INPUT_191       => INPUT_191,
    INPUT_192       => INPUT_192,
    INPUT_193       => INPUT_193,
    INPUT_194       => INPUT_194,
    INPUT_195       => INPUT_195,
    INPUT_196       => INPUT_196,
    INPUT_197       => INPUT_197,
    INPUT_198       => INPUT_198,
    INPUT_199       => INPUT_199,
    INPUT_200       => INPUT_200,
    INPUT_201       => INPUT_201,
    INPUT_202       => INPUT_202,
    INPUT_203       => INPUT_203,
    INPUT_204       => INPUT_204,
    INPUT_205       => INPUT_205,
    INPUT_206       => INPUT_206,
    INPUT_207       => INPUT_207,
    INPUT_208       => INPUT_208,
    INPUT_209       => INPUT_209,
    INPUT_210       => INPUT_210,
    INPUT_211       => INPUT_211,
    INPUT_212       => INPUT_212,
    INPUT_213       => INPUT_213,
    INPUT_214       => INPUT_214,
    INPUT_215       => INPUT_215,
    INPUT_216       => INPUT_216,
    INPUT_217       => INPUT_217,
    INPUT_218       => INPUT_218,
    INPUT_219       => INPUT_219,
    INPUT_220       => INPUT_220,
    INPUT_221       => INPUT_221,
    INPUT_222       => INPUT_222,
    INPUT_223       => INPUT_223,
    INPUT_224       => INPUT_224,
    INPUT_225       => INPUT_225,
    INPUT_226       => INPUT_226,
    INPUT_227       => INPUT_227,
    INPUT_228       => INPUT_228,
    INPUT_229       => INPUT_229,
    INPUT_230       => INPUT_230,
    INPUT_231       => INPUT_231,
    INPUT_232       => INPUT_232,
    INPUT_233       => INPUT_233,
    INPUT_234       => INPUT_234,
    INPUT_235       => INPUT_235,
    INPUT_236       => INPUT_236,
    INPUT_237       => INPUT_237,
    INPUT_238       => INPUT_238,
    INPUT_239       => INPUT_239,
    INPUT_240       => INPUT_240,
    INPUT_241       => INPUT_241,
    INPUT_242       => INPUT_242,
    INPUT_243       => INPUT_243,
    INPUT_244       => INPUT_244,
    INPUT_245       => INPUT_245,
    INPUT_246       => INPUT_246,
    INPUT_247       => INPUT_247,
    INPUT_248       => INPUT_248,
    INPUT_249       => INPUT_249,
    INPUT_250       => INPUT_250,
    INPUT_251       => INPUT_251,
    INPUT_252       => INPUT_252,
    INPUT_253       => INPUT_253,
    INPUT_254       => INPUT_254,
    INPUT_255       => INPUT_255,
    INPUT_256       => INPUT_256,
    INPUT_257       => INPUT_257,
    INPUT_258       => INPUT_258,
    INPUT_259       => INPUT_259,
    INPUT_260       => INPUT_260,
    INPUT_261       => INPUT_261,
    INPUT_262       => INPUT_262,
    INPUT_263       => INPUT_263,
    INPUT_264       => INPUT_264,
    INPUT_265       => INPUT_265,
    INPUT_266       => INPUT_266,
    INPUT_267       => INPUT_267,
    INPUT_268       => INPUT_268,
    INPUT_269       => INPUT_269,
    INPUT_270       => INPUT_270,
    INPUT_271       => INPUT_271,
    INPUT_272       => INPUT_272,
    INPUT_273       => INPUT_273,
    INPUT_274       => INPUT_274,
    INPUT_275       => INPUT_275,
    INPUT_276       => INPUT_276,
    INPUT_277       => INPUT_277,
    INPUT_278       => INPUT_278,
    INPUT_279       => INPUT_279,
    INPUT_280       => INPUT_280,
    INPUT_281       => INPUT_281,
    INPUT_282       => INPUT_282,
    INPUT_283       => INPUT_283,
    INPUT_284       => INPUT_284,
    INPUT_285       => INPUT_285,
    INPUT_286       => INPUT_286,
    INPUT_287       => INPUT_287,
    INPUT_288       => INPUT_288,
    INPUT_289       => INPUT_289,
    INPUT_290       => INPUT_290,
    INPUT_291       => INPUT_291,
    INPUT_292       => INPUT_292,
    INPUT_293       => INPUT_293,
    INPUT_294       => INPUT_294,
    INPUT_295       => INPUT_295,
    INPUT_296       => INPUT_296,
    INPUT_297       => INPUT_297,
    INPUT_298       => INPUT_298,
    INPUT_299       => INPUT_299,
    INPUT_300       => INPUT_300,
    INPUT_301       => INPUT_301,
    INPUT_302       => INPUT_302,
    INPUT_303       => INPUT_303,
    INPUT_304       => INPUT_304,
    INPUT_305       => INPUT_305,
    INPUT_306       => INPUT_306,
    INPUT_307       => INPUT_307,
    INPUT_308       => INPUT_308,
    INPUT_309       => INPUT_309,
    INPUT_310       => INPUT_310,
    INPUT_311       => INPUT_311,
    INPUT_312       => INPUT_312,
    INPUT_313       => INPUT_313,
    INPUT_314       => INPUT_314,
    INPUT_315       => INPUT_315,
    INPUT_316       => INPUT_316,
    INPUT_317       => INPUT_317,
    INPUT_318       => INPUT_318,
    INPUT_319       => INPUT_319,
    INPUT_320       => INPUT_320,
    INPUT_321       => INPUT_321,
    INPUT_322       => INPUT_322,
    INPUT_323       => INPUT_323,
    INPUT_324       => INPUT_324,
    INPUT_325       => INPUT_325,
    INPUT_326       => INPUT_326,
    INPUT_327       => INPUT_327,
    INPUT_328       => INPUT_328,
    INPUT_329       => INPUT_329,
    INPUT_330       => INPUT_330,
    INPUT_331       => INPUT_331,
    INPUT_332       => INPUT_332,
    INPUT_333       => INPUT_333,
    INPUT_334       => INPUT_334,
    INPUT_335       => INPUT_335,
    INPUT_336       => INPUT_336,
    INPUT_337       => INPUT_337,
    INPUT_338       => INPUT_338,
    INPUT_339       => INPUT_339,
    INPUT_340       => INPUT_340,
    INPUT_341       => INPUT_341,
    INPUT_342       => INPUT_342,
    INPUT_343       => INPUT_343,
    INPUT_344       => INPUT_344,
    INPUT_345       => INPUT_345,
    INPUT_346       => INPUT_346,
    INPUT_347       => INPUT_347,
    INPUT_348       => INPUT_348,
    INPUT_349       => INPUT_349,
    INPUT_350       => INPUT_350,
    INPUT_351       => INPUT_351,
    INPUT_352       => INPUT_352,
    INPUT_353       => INPUT_353,
    INPUT_354       => INPUT_354,
    INPUT_355       => INPUT_355,
    INPUT_356       => INPUT_356,
    INPUT_357       => INPUT_357,
    INPUT_358       => INPUT_358,
    INPUT_359       => INPUT_359,
    INPUT_360       => INPUT_360,
    INPUT_361       => INPUT_361,
    INPUT_362       => INPUT_362,
    INPUT_363       => INPUT_363,
    INPUT_364       => INPUT_364,
    INPUT_365       => INPUT_365,
    INPUT_366       => INPUT_366,
    INPUT_367       => INPUT_367,
    INPUT_368       => INPUT_368,
    INPUT_369       => INPUT_369,
    INPUT_370       => INPUT_370,
    INPUT_371       => INPUT_371,
    INPUT_372       => INPUT_372,
    INPUT_373       => INPUT_373,
    INPUT_374       => INPUT_374,
    INPUT_375       => INPUT_375,
    INPUT_376       => INPUT_376,
    INPUT_377       => INPUT_377,
    INPUT_378       => INPUT_378,
    INPUT_379       => INPUT_379,
    INPUT_380       => INPUT_380,
    INPUT_381       => INPUT_381,
    INPUT_382       => INPUT_382,
    INPUT_383       => INPUT_383,
    INPUT_384       => INPUT_384,
    INPUT_385       => INPUT_385,
    INPUT_386       => INPUT_386,
    INPUT_387       => INPUT_387,
    INPUT_388       => INPUT_388,
    INPUT_389       => INPUT_389,
    INPUT_390       => INPUT_390,
    INPUT_391       => INPUT_391,
    INPUT_392       => INPUT_392,
    INPUT_393       => INPUT_393,
    INPUT_394       => INPUT_394,
    INPUT_395       => INPUT_395,
    INPUT_396       => INPUT_396,
    INPUT_397       => INPUT_397,
    INPUT_398       => INPUT_398,
    INPUT_399       => INPUT_399,
    INPUT_400       => INPUT_400,
    INPUT_401       => INPUT_401,
    INPUT_402       => INPUT_402,
    INPUT_403       => INPUT_403,
    INPUT_404       => INPUT_404,
    INPUT_405       => INPUT_405,
    INPUT_406       => INPUT_406,
    INPUT_407       => INPUT_407,
    INPUT_408       => INPUT_408,
    INPUT_409       => INPUT_409,
    INPUT_410       => INPUT_410,
    INPUT_411       => INPUT_411,
    INPUT_412       => INPUT_412,
    INPUT_413       => INPUT_413,
    INPUT_414       => INPUT_414,
    INPUT_415       => INPUT_415,
    INPUT_416       => INPUT_416,
    INPUT_417       => INPUT_417,
    INPUT_418       => INPUT_418,
    INPUT_419       => INPUT_419,
    INPUT_420       => INPUT_420,
    INPUT_421       => INPUT_421,
    INPUT_422       => INPUT_422,
    INPUT_423       => INPUT_423,
    INPUT_424       => INPUT_424,
    INPUT_425       => INPUT_425,
    INPUT_426       => INPUT_426,
    INPUT_427       => INPUT_427,
    INPUT_428       => INPUT_428,
    INPUT_429       => INPUT_429,
    INPUT_430       => INPUT_430,
    INPUT_431       => INPUT_431,
    INPUT_432       => INPUT_432,
    INPUT_433       => INPUT_433,
    INPUT_434       => INPUT_434,
    INPUT_435       => INPUT_435,
    INPUT_436       => INPUT_436,
    INPUT_437       => INPUT_437,
    INPUT_438       => INPUT_438,
    INPUT_439       => INPUT_439,
    INPUT_440       => INPUT_440,
    INPUT_441       => INPUT_441,
    INPUT_442       => INPUT_442,
    INPUT_443       => INPUT_443,
    INPUT_444       => INPUT_444,
    INPUT_445       => INPUT_445,
    INPUT_446       => INPUT_446,
    INPUT_447       => INPUT_447,
    INPUT_448       => INPUT_448,
    INPUT_449       => INPUT_449,
    INPUT_450       => INPUT_450,
    INPUT_451       => INPUT_451,
    INPUT_452       => INPUT_452,
    INPUT_453       => INPUT_453,
    INPUT_454       => INPUT_454,
    INPUT_455       => INPUT_455,
    INPUT_456       => INPUT_456,
    INPUT_457       => INPUT_457,
    INPUT_458       => INPUT_458,
    INPUT_459       => INPUT_459,
    INPUT_460       => INPUT_460,
    INPUT_461       => INPUT_461,
    INPUT_462       => INPUT_462,
    INPUT_463       => INPUT_463,
    INPUT_464       => INPUT_464,
    INPUT_465       => INPUT_465,
    INPUT_466       => INPUT_466,
    INPUT_467       => INPUT_467,
    INPUT_468       => INPUT_468,
    INPUT_469       => INPUT_469,
    INPUT_470       => INPUT_470,
    INPUT_471       => INPUT_471,
    INPUT_472       => INPUT_472,
    INPUT_473       => INPUT_473,
    INPUT_474       => INPUT_474,
    INPUT_475       => INPUT_475,
    INPUT_476       => INPUT_476,
    INPUT_477       => INPUT_477,
    INPUT_478       => INPUT_478,
    INPUT_479       => INPUT_479,
    INPUT_480       => INPUT_480,
    INPUT_481       => INPUT_481,
    INPUT_482       => INPUT_482,
    INPUT_483       => INPUT_483,
    INPUT_484       => INPUT_484,
    INPUT_485       => INPUT_485,
    INPUT_486       => INPUT_486,
    INPUT_487       => INPUT_487,
    INPUT_488       => INPUT_488,
    INPUT_489       => INPUT_489,
    INPUT_490       => INPUT_490,
    INPUT_491       => INPUT_491,
    INPUT_492       => INPUT_492,
    INPUT_493       => INPUT_493,
    INPUT_494       => INPUT_494,
    INPUT_495       => INPUT_495,
    INPUT_496       => INPUT_496,
    INPUT_497       => INPUT_497,
    INPUT_498       => INPUT_498,
    INPUT_499       => INPUT_499,
    INPUT_500       => INPUT_500,
    INPUT_501       => INPUT_501,
    INPUT_502       => INPUT_502,
    INPUT_503       => INPUT_503,
    INPUT_504       => INPUT_504,
    INPUT_505       => INPUT_505,
    INPUT_506       => INPUT_506,
    INPUT_507       => INPUT_507,
    INPUT_508       => INPUT_508,
    INPUT_509       => INPUT_509,
    INPUT_510       => INPUT_510,
    INPUT_511       => INPUT_511,
    INPUT_512       => INPUT_512,
    INPUT_513       => INPUT_513,
    INPUT_514       => INPUT_514,
    INPUT_515       => INPUT_515,
    INPUT_516       => INPUT_516,
    INPUT_517       => INPUT_517,
    INPUT_518       => INPUT_518,
    INPUT_519       => INPUT_519,
    INPUT_520       => INPUT_520,
    INPUT_521       => INPUT_521,
    INPUT_522       => INPUT_522,
    INPUT_523       => INPUT_523,
    INPUT_524       => INPUT_524,
    INPUT_525       => INPUT_525,
    INPUT_526       => INPUT_526,
    INPUT_527       => INPUT_527,
    INPUT_528       => INPUT_528,
    INPUT_529       => INPUT_529,
    INPUT_530       => INPUT_530,
    INPUT_531       => INPUT_531,
    INPUT_532       => INPUT_532,
    INPUT_533       => INPUT_533,
    INPUT_534       => INPUT_534,
    INPUT_535       => INPUT_535,
    INPUT_536       => INPUT_536,
    INPUT_537       => INPUT_537,
    INPUT_538       => INPUT_538,
    INPUT_539       => INPUT_539,
    INPUT_540       => INPUT_540,
    INPUT_541       => INPUT_541,
    INPUT_542       => INPUT_542,
    INPUT_543       => INPUT_543,
    INPUT_544       => INPUT_544,
    INPUT_545       => INPUT_545,
    INPUT_546       => INPUT_546,
    INPUT_547       => INPUT_547,
    INPUT_548       => INPUT_548,
    INPUT_549       => INPUT_549,
    INPUT_550       => INPUT_550,
    INPUT_551       => INPUT_551,
    INPUT_552       => INPUT_552,
    INPUT_553       => INPUT_553,
    INPUT_554       => INPUT_554,
    INPUT_555       => INPUT_555,
    INPUT_556       => INPUT_556,
    INPUT_557       => INPUT_557,
    INPUT_558       => INPUT_558,
    INPUT_559       => INPUT_559,
    INPUT_560       => INPUT_560,
    INPUT_561       => INPUT_561,
    INPUT_562       => INPUT_562,
    INPUT_563       => INPUT_563,
    INPUT_564       => INPUT_564,
    INPUT_565       => INPUT_565,
    INPUT_566       => INPUT_566,
    INPUT_567       => INPUT_567,
    INPUT_568       => INPUT_568,
    INPUT_569       => INPUT_569,
    INPUT_570       => INPUT_570,
    INPUT_571       => INPUT_571,
    INPUT_572       => INPUT_572,
    INPUT_573       => INPUT_573,
    INPUT_574       => INPUT_574,
    INPUT_575       => INPUT_575,
    INPUT_576       => INPUT_576,
    INPUT_577       => INPUT_577,
    INPUT_578       => INPUT_578,
    INPUT_579       => INPUT_579,
    INPUT_580       => INPUT_580,
    INPUT_581       => INPUT_581,
    INPUT_582       => INPUT_582,
    INPUT_583       => INPUT_583,
    INPUT_584       => INPUT_584,
    INPUT_585       => INPUT_585,
    INPUT_586       => INPUT_586,
    INPUT_587       => INPUT_587,
    INPUT_588       => INPUT_588,
    INPUT_589       => INPUT_589,
    INPUT_590       => INPUT_590,
    INPUT_591       => INPUT_591,
    INPUT_592       => INPUT_592,
    INPUT_593       => INPUT_593,
    INPUT_594       => INPUT_594,
    INPUT_595       => INPUT_595,
    INPUT_596       => INPUT_596,
    INPUT_597       => INPUT_597,
    INPUT_598       => INPUT_598,
    INPUT_599       => INPUT_599,
    INPUT_600       => INPUT_600,
    INPUT_601       => INPUT_601,
    INPUT_602       => INPUT_602,
    INPUT_603       => INPUT_603,
    INPUT_604       => INPUT_604,
    INPUT_605       => INPUT_605,
    INPUT_606       => INPUT_606,
    INPUT_607       => INPUT_607,
    INPUT_608       => INPUT_608,
    INPUT_609       => INPUT_609,
    INPUT_610       => INPUT_610,
    INPUT_611       => INPUT_611,
    INPUT_612       => INPUT_612,
    INPUT_613       => INPUT_613,
    INPUT_614       => INPUT_614,
    INPUT_615       => INPUT_615,
    INPUT_616       => INPUT_616,
    INPUT_617       => INPUT_617,
    INPUT_618       => INPUT_618,
    INPUT_619       => INPUT_619,
    INPUT_620       => INPUT_620,
    INPUT_621       => INPUT_621,
    INPUT_622       => INPUT_622,
    INPUT_623       => INPUT_623,
    INPUT_624       => INPUT_624,
    INPUT_625       => INPUT_625,
    INPUT_626       => INPUT_626,
    INPUT_627       => INPUT_627,
    INPUT_628       => INPUT_628,
    INPUT_629       => INPUT_629,
    INPUT_630       => INPUT_630,
    INPUT_631       => INPUT_631,
    INPUT_632       => INPUT_632,
    INPUT_633       => INPUT_633,
    INPUT_634       => INPUT_634,
    INPUT_635       => INPUT_635,
    INPUT_636       => INPUT_636,
    INPUT_637       => INPUT_637,
    INPUT_638       => INPUT_638,
    INPUT_639       => INPUT_639,
    INPUT_640       => INPUT_640,
    INPUT_641       => INPUT_641,
    INPUT_642       => INPUT_642,
    INPUT_643       => INPUT_643,
    INPUT_644       => INPUT_644,
    INPUT_645       => INPUT_645,
    INPUT_646       => INPUT_646,
    INPUT_647       => INPUT_647,
    INPUT_648       => INPUT_648,
    INPUT_649       => INPUT_649,
    INPUT_650       => INPUT_650,
    INPUT_651       => INPUT_651,
    INPUT_652       => INPUT_652,
    INPUT_653       => INPUT_653,
    INPUT_654       => INPUT_654,
    OUTPUT      => OUTPUT,
    OUTPUT_2 => OUTPUT_2,
    VALID     => VALID,
    START     => START,
    RUNTIME     => RUNTIME,
    FINISHED    => FINISHED,
    BUSY      => BUSY,
    OUTPUT_CYCLE  => OUTPUT_CYCLE
  );
  
Clk_gen : PROCESS
BEGIN
  SYS_CLK <= '1';
  WAIT FOR clk_per/2;
  SYS_CLK <= '0';
  WAIT FOR clk_per/2;
END PROCESS;

Rst_gen : PROCESS
BEGIN
  SYS_RST <= '1';
  WAIT UNTIL rising_edge(SYS_CLK);
  SYS_RST <= '0';
  WAIT;
END PROCESS;  


tb : PROCESS

   file output_x : TEXT open WRITE_MODE is "x.out";
   file output_lpr : TEXT open WRITE_MODE is "LPR.out";
   variable output_line: line;

BEGIN
  --Initialisation of input signals
  steps <= INPUT_1;
  runs <= INPUT_2;

  BUSY <= '0';
  
  toggle_start(SYS_CLK, START);

  while i < to_integer(unsigned(RUNS))*CHAINS loop
    if VALID = '1' then
      i <= i +1;
      hwrite(output_line, OUTPUT);
      writeline(output_x, output_line);
      hwrite(output_line, OUTPUT_2);
      writeline(output_x, output_line);
    end if;
    wait for clk_per;
  end loop ; 

  i <= 0;
  
  while i < (to_integer(unsigned(STEPS))/BLOCKS)*to_integer(unsigned(RUNS))*CHAINS*BLOCKS loop
    if VALID = '1' then
      i <= i +1;
      hwrite(output_line, OUTPUT);
      writeline(output_lpr, output_line);
      hwrite(output_line, OUTPUT_2);
      writeline(output_lpr, output_line);
    end if;
    wait for clk_per;
  end loop ;

  WAIT UNTIL rising_edge(FINISHED);
  -- wait_for(SYS_CLK,5);
  
  -- --BUSY signal test
  
  -- BUSY <= '1';
  
  -- toggle_start(SYS_CLK, START);
  -- wait_for(SYS_CLK,20);
  
  -- BUSY <= '0';
  
  -- WAIT UNTIL rising_edge(FINISHED);
  -- wait_for(SYS_CLK,5);
  
  REPORT "TEST FINISHED." SEVERITY failure;
END PROCESS;

END ARCHITECTURE test_bench;