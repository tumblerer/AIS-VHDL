library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Beta_pack is
	
	type beta_type is array (0 downto 20) of std_logic_vector(63 downto 0);

	constant 
end package ; -- Beta 