--------------------------------------------------------------------------------
--                               Compressor_2_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_2_2 is
   port ( X0 : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_2_2 is
signal X :  std_logic_vector(1 downto 0);
begin
   X <=X0 ;
   with X select R <= 
      "00" when "00", 
      "01" when "01", 
      "01" when "10", 
      "10" when "11", 
      "--" when others;

end architecture;

--------------------------------------------------------------------------------
--                               Compressor_3_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2 is
   port ( X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2 is
signal X :  std_logic_vector(2 downto 0);
begin
   X <=X0 ;
   with X select R <= 
      "00" when "000", 
      "01" when "001", 
      "01" when "010", 
      "10" when "011", 
      "01" when "100", 
      "10" when "101", 
      "10" when "110", 
      "11" when "111", 
      "--" when others;

end architecture;

--------------------------------------------------------------------------------
--                               LZOC_52_6_uid3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_52_6_uid3 is
   port ( clk, rst : in std_logic;
          I : in  std_logic_vector(51 downto 0);
          OZB : in std_logic;
          O : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of LZOC_52_6_uid3 is
signal sozb, sozb_d1, sozb_d2, sozb_d3 : std_logic;
signal level6 :  std_logic_vector(63 downto 0);
signal digit6, digit6_d1, digit6_d2, digit6_d3 : std_logic;
signal level5, level5_d1 :  std_logic_vector(31 downto 0);
signal digit5, digit5_d1, digit5_d2 : std_logic;
signal level4, level4_d1 :  std_logic_vector(15 downto 0);
signal digit4, digit4_d1, digit4_d2 : std_logic;
signal level3 :  std_logic_vector(7 downto 0);
signal digit3, digit3_d1 : std_logic;
signal level2 :  std_logic_vector(3 downto 0);
signal digit2, digit2_d1 : std_logic;
signal level1, level1_d1 :  std_logic_vector(1 downto 0);
signal digit1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sozb_d1 <=  sozb;
            sozb_d2 <=  sozb_d1;
            sozb_d3 <=  sozb_d2;
            digit6_d1 <=  digit6;
            digit6_d2 <=  digit6_d1;
            digit6_d3 <=  digit6_d2;
            level5_d1 <=  level5;
            digit5_d1 <=  digit5;
            digit5_d2 <=  digit5_d1;
            level4_d1 <=  level4;
            digit4_d1 <=  digit4;
            digit4_d2 <=  digit4_d1;
            digit3_d1 <=  digit3;
            digit2_d1 <=  digit2;
            level1_d1 <=  level1;
         end if;
      end process;
   sozb <= OZB;
   level6<= I& (11 downto 0 => not(sozb));
   digit6<= '1' when level6(63 downto 32) = (63 downto 32 => sozb) else '0';
   level5<= level6(31 downto 0) when digit6='1' else level6(63 downto 32);
   ----------------Synchro barrier, entering cycle 1----------------
   digit5<= '1' when level5_d1(31 downto 16) = (31 downto 16 => sozb_d1) else '0';
   level4<= level5_d1(15 downto 0) when digit5='1' else level5_d1(31 downto 16);
   digit4<= '1' when level4(15 downto 8) = (15 downto 8 => sozb_d1) else '0';
   ----------------Synchro barrier, entering cycle 2----------------
   level3<= level4_d1(7 downto 0) when digit4_d1='1' else level4_d1(15 downto 8);
   digit3<= '1' when level3(7 downto 4) = (7 downto 4 => sozb_d2) else '0';
   level2<= level3(3 downto 0) when digit3='1' else level3(7 downto 4);
   digit2<= '1' when level2(3 downto 2) = (3 downto 2 => sozb_d2) else '0';
   level1<= level2(1 downto 0) when digit2='1' else level2(3 downto 2);
   ----------------Synchro barrier, entering cycle 3----------------
   digit1<= '1' when level1_d1(1 downto 1) = (1 downto 1 => sozb_d3) else '0';
   O <= digit6_d3 & digit5_d2 & digit4_d2 & digit3_d1 & digit2_d1 & digit1;
end architecture;

--------------------------------------------------------------------------------
--                       LeftShifter_27_by_max_27_uid6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter_27_by_max_27_uid6 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(26 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(53 downto 0)   );
end entity;

architecture arch of LeftShifter_27_by_max_27_uid6 is
signal level0, level0_d1 :  std_logic_vector(26 downto 0);
signal ps, ps_d1 :  std_logic_vector(4 downto 0);
signal level1 :  std_logic_vector(27 downto 0);
signal level2 :  std_logic_vector(29 downto 0);
signal level3 :  std_logic_vector(33 downto 0);
signal level4 :  std_logic_vector(41 downto 0);
signal level5 :  std_logic_vector(57 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            level0_d1 <=  level0;
            ps_d1 <=  ps;
         end if;
      end process;
   level0<= X;
   ps<= S;
   ----------------Synchro barrier, entering cycle 1----------------
   level1<= level0_d1 & (0 downto 0 => '0') when ps_d1(0)= '1' else     (0 downto 0 => '0') & level0_d1;
   level2<= level1 & (1 downto 0 => '0') when ps_d1(1)= '1' else     (1 downto 0 => '0') & level1;
   level3<= level2 & (3 downto 0 => '0') when ps_d1(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3;
   level5<= level4 & (15 downto 0 => '0') when ps_d1(4)= '1' else     (15 downto 0 => '0') & level4;
   R <= level5(53 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                              InvTable_0_11_12
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity InvTable_0_11_12 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          Y : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of InvTable_0_11_12 is
   -- Build a 2-D array type for the RoM
   subtype word_t is std_logic_vector(11 downto 0);
   type memory_t is array(0 to 2047) of word_t;
   function init_rom
      return memory_t is 
      variable tmp : memory_t := (
   "100000000000",
   "100000000000",
   "011111111111",
   "011111111110",
   "011111111101",
   "011111111100",
   "011111111011",
   "011111111010",
   "011111111001",
   "011111111000",
   "011111110111",
   "011111110110",
   "011111110101",
   "011111110100",
   "011111110011",
   "011111110010",
   "011111110001",
   "011111110000",
   "011111101111",
   "011111101110",
   "011111101101",
   "011111101100",
   "011111101011",
   "011111101010",
   "011111101001",
   "011111101000",
   "011111100111",
   "011111100110",
   "011111100101",
   "011111100100",
   "011111100011",
   "011111100010",
   "011111100001",
   "011111100000",
   "011111011111",
   "011111011110",
   "011111011101",
   "011111011100",
   "011111011011",
   "011111011010",
   "011111011001",
   "011111011000",
   "011111010111",
   "011111010110",
   "011111010101",
   "011111010100",
   "011111010100",
   "011111010011",
   "011111010010",
   "011111010001",
   "011111010000",
   "011111001111",
   "011111001110",
   "011111001101",
   "011111001100",
   "011111001011",
   "011111001010",
   "011111001001",
   "011111001000",
   "011111000111",
   "011111000110",
   "011111000101",
   "011111000100",
   "011111000011",
   "011111000010",
   "011111000001",
   "011111000001",
   "011111000000",
   "011110111111",
   "011110111110",
   "011110111101",
   "011110111100",
   "011110111011",
   "011110111010",
   "011110111001",
   "011110111000",
   "011110110111",
   "011110110110",
   "011110110101",
   "011110110100",
   "011110110100",
   "011110110011",
   "011110110010",
   "011110110001",
   "011110110000",
   "011110101111",
   "011110101110",
   "011110101101",
   "011110101100",
   "011110101011",
   "011110101010",
   "011110101001",
   "011110101000",
   "011110101000",
   "011110100111",
   "011110100110",
   "011110100101",
   "011110100100",
   "011110100011",
   "011110100010",
   "011110100001",
   "011110100000",
   "011110011111",
   "011110011110",
   "011110011110",
   "011110011101",
   "011110011100",
   "011110011011",
   "011110011010",
   "011110011001",
   "011110011000",
   "011110010111",
   "011110010110",
   "011110010101",
   "011110010101",
   "011110010100",
   "011110010011",
   "011110010010",
   "011110010001",
   "011110010000",
   "011110001111",
   "011110001110",
   "011110001101",
   "011110001100",
   "011110001100",
   "011110001011",
   "011110001010",
   "011110001001",
   "011110001000",
   "011110000111",
   "011110000110",
   "011110000101",
   "011110000100",
   "011110000100",
   "011110000011",
   "011110000010",
   "011110000001",
   "011110000000",
   "011101111111",
   "011101111110",
   "011101111101",
   "011101111101",
   "011101111100",
   "011101111011",
   "011101111010",
   "011101111001",
   "011101111000",
   "011101110111",
   "011101110110",
   "011101110110",
   "011101110101",
   "011101110100",
   "011101110011",
   "011101110010",
   "011101110001",
   "011101110000",
   "011101110000",
   "011101101111",
   "011101101110",
   "011101101101",
   "011101101100",
   "011101101011",
   "011101101010",
   "011101101010",
   "011101101001",
   "011101101000",
   "011101100111",
   "011101100110",
   "011101100101",
   "011101100100",
   "011101100100",
   "011101100011",
   "011101100010",
   "011101100001",
   "011101100000",
   "011101011111",
   "011101011110",
   "011101011110",
   "011101011101",
   "011101011100",
   "011101011011",
   "011101011010",
   "011101011001",
   "011101011001",
   "011101011000",
   "011101010111",
   "011101010110",
   "011101010101",
   "011101010100",
   "011101010011",
   "011101010011",
   "011101010010",
   "011101010001",
   "011101010000",
   "011101001111",
   "011101001110",
   "011101001110",
   "011101001101",
   "011101001100",
   "011101001011",
   "011101001010",
   "011101001001",
   "011101001001",
   "011101001000",
   "011101000111",
   "011101000110",
   "011101000101",
   "011101000101",
   "011101000100",
   "011101000011",
   "011101000010",
   "011101000001",
   "011101000000",
   "011101000000",
   "011100111111",
   "011100111110",
   "011100111101",
   "011100111100",
   "011100111011",
   "011100111011",
   "011100111010",
   "011100111001",
   "011100111000",
   "011100110111",
   "011100110111",
   "011100110110",
   "011100110101",
   "011100110100",
   "011100110011",
   "011100110011",
   "011100110010",
   "011100110001",
   "011100110000",
   "011100101111",
   "011100101110",
   "011100101110",
   "011100101101",
   "011100101100",
   "011100101011",
   "011100101010",
   "011100101010",
   "011100101001",
   "011100101000",
   "011100100111",
   "011100100110",
   "011100100110",
   "011100100101",
   "011100100100",
   "011100100011",
   "011100100010",
   "011100100010",
   "011100100001",
   "011100100000",
   "011100011111",
   "011100011111",
   "011100011110",
   "011100011101",
   "011100011100",
   "011100011011",
   "011100011011",
   "011100011010",
   "011100011001",
   "011100011000",
   "011100010111",
   "011100010111",
   "011100010110",
   "011100010101",
   "011100010100",
   "011100010100",
   "011100010011",
   "011100010010",
   "011100010001",
   "011100010000",
   "011100010000",
   "011100001111",
   "011100001110",
   "011100001101",
   "011100001101",
   "011100001100",
   "011100001011",
   "011100001010",
   "011100001001",
   "011100001001",
   "011100001000",
   "011100000111",
   "011100000110",
   "011100000110",
   "011100000101",
   "011100000100",
   "011100000011",
   "011100000010",
   "011100000010",
   "011100000001",
   "011100000000",
   "011011111111",
   "011011111111",
   "011011111110",
   "011011111101",
   "011011111100",
   "011011111100",
   "011011111011",
   "011011111010",
   "011011111001",
   "011011111001",
   "011011111000",
   "011011110111",
   "011011110110",
   "011011110110",
   "011011110101",
   "011011110100",
   "011011110011",
   "011011110011",
   "011011110010",
   "011011110001",
   "011011110000",
   "011011101111",
   "011011101111",
   "011011101110",
   "011011101101",
   "011011101100",
   "011011101100",
   "011011101011",
   "011011101010",
   "011011101010",
   "011011101001",
   "011011101000",
   "011011100111",
   "011011100111",
   "011011100110",
   "011011100101",
   "011011100100",
   "011011100100",
   "011011100011",
   "011011100010",
   "011011100001",
   "011011100001",
   "011011100000",
   "011011011111",
   "011011011110",
   "011011011110",
   "011011011101",
   "011011011100",
   "011011011011",
   "011011011011",
   "011011011010",
   "011011011001",
   "011011011001",
   "011011011000",
   "011011010111",
   "011011010110",
   "011011010110",
   "011011010101",
   "011011010100",
   "011011010011",
   "011011010011",
   "011011010010",
   "011011010001",
   "011011010000",
   "011011010000",
   "011011001111",
   "011011001110",
   "011011001110",
   "011011001101",
   "011011001100",
   "011011001011",
   "011011001011",
   "011011001010",
   "011011001001",
   "011011001001",
   "011011001000",
   "011011000111",
   "011011000110",
   "011011000110",
   "011011000101",
   "011011000100",
   "011011000100",
   "011011000011",
   "011011000010",
   "011011000001",
   "011011000001",
   "011011000000",
   "011010111111",
   "011010111111",
   "011010111110",
   "011010111101",
   "011010111100",
   "011010111100",
   "011010111011",
   "011010111010",
   "011010111010",
   "011010111001",
   "011010111000",
   "011010110111",
   "011010110111",
   "011010110110",
   "011010110101",
   "011010110101",
   "011010110100",
   "011010110011",
   "011010110011",
   "011010110010",
   "011010110001",
   "011010110000",
   "011010110000",
   "011010101111",
   "011010101110",
   "011010101110",
   "011010101101",
   "011010101100",
   "011010101100",
   "011010101011",
   "011010101010",
   "011010101010",
   "011010101001",
   "011010101000",
   "011010100111",
   "011010100111",
   "011010100110",
   "011010100101",
   "011010100101",
   "011010100100",
   "011010100011",
   "011010100011",
   "011010100010",
   "011010100001",
   "011010100001",
   "011010100000",
   "011010011111",
   "011010011110",
   "011010011110",
   "011010011101",
   "011010011100",
   "011010011100",
   "011010011011",
   "011010011010",
   "011010011010",
   "011010011001",
   "011010011000",
   "011010011000",
   "011010010111",
   "011010010110",
   "011010010110",
   "011010010101",
   "011010010100",
   "011010010100",
   "011010010011",
   "011010010010",
   "011010010010",
   "011010010001",
   "011010010000",
   "011010010000",
   "011010001111",
   "011010001110",
   "011010001110",
   "011010001101",
   "011010001100",
   "011010001100",
   "011010001011",
   "011010001010",
   "011010001010",
   "011010001001",
   "011010001000",
   "011010001000",
   "011010000111",
   "011010000110",
   "011010000110",
   "011010000101",
   "011010000100",
   "011010000100",
   "011010000011",
   "011010000010",
   "011010000010",
   "011010000001",
   "011010000000",
   "011010000000",
   "011001111111",
   "011001111110",
   "011001111110",
   "011001111101",
   "011001111100",
   "011001111100",
   "011001111011",
   "011001111010",
   "011001111010",
   "011001111001",
   "011001111000",
   "011001111000",
   "011001110111",
   "011001110110",
   "011001110110",
   "011001110101",
   "011001110100",
   "011001110100",
   "011001110011",
   "011001110011",
   "011001110010",
   "011001110001",
   "011001110001",
   "011001110000",
   "011001101111",
   "011001101111",
   "011001101110",
   "011001101101",
   "011001101101",
   "011001101100",
   "011001101011",
   "011001101011",
   "011001101010",
   "011001101001",
   "011001101001",
   "011001101000",
   "011001101000",
   "011001100111",
   "011001100110",
   "011001100110",
   "011001100101",
   "011001100100",
   "011001100100",
   "011001100011",
   "011001100010",
   "011001100010",
   "011001100001",
   "011001100001",
   "011001100000",
   "011001011111",
   "011001011111",
   "011001011110",
   "011001011101",
   "011001011101",
   "011001011100",
   "011001011011",
   "011001011011",
   "011001011010",
   "011001011010",
   "011001011001",
   "011001011000",
   "011001011000",
   "011001010111",
   "011001010110",
   "011001010110",
   "011001010101",
   "011001010101",
   "011001010100",
   "011001010011",
   "011001010011",
   "011001010010",
   "011001010001",
   "011001010001",
   "011001010000",
   "011001010000",
   "011001001111",
   "011001001110",
   "011001001110",
   "011001001101",
   "011001001100",
   "011001001100",
   "011001001011",
   "011001001011",
   "011001001010",
   "011001001001",
   "011001001001",
   "011001001000",
   "011001001000",
   "011001000111",
   "011001000110",
   "011001000110",
   "011001000101",
   "011001000100",
   "011001000100",
   "011001000011",
   "011001000011",
   "011001000010",
   "011001000001",
   "011001000001",
   "011001000000",
   "011001000000",
   "011000111111",
   "011000111110",
   "011000111110",
   "011000111101",
   "011000111101",
   "011000111100",
   "011000111011",
   "011000111011",
   "011000111010",
   "011000111001",
   "011000111001",
   "011000111000",
   "011000111000",
   "011000110111",
   "011000110110",
   "011000110110",
   "011000110101",
   "011000110101",
   "011000110100",
   "011000110011",
   "011000110011",
   "011000110010",
   "011000110010",
   "011000110001",
   "011000110000",
   "011000110000",
   "011000101111",
   "011000101111",
   "011000101110",
   "011000101101",
   "011000101101",
   "011000101100",
   "011000101100",
   "011000101011",
   "011000101010",
   "011000101010",
   "011000101001",
   "011000101001",
   "011000101000",
   "011000101000",
   "011000100111",
   "011000100110",
   "011000100110",
   "011000100101",
   "011000100101",
   "011000100100",
   "011000100011",
   "011000100011",
   "011000100010",
   "011000100010",
   "011000100001",
   "011000100000",
   "011000100000",
   "011000011111",
   "011000011111",
   "011000011110",
   "011000011110",
   "011000011101",
   "011000011100",
   "011000011100",
   "011000011011",
   "011000011011",
   "011000011010",
   "011000011001",
   "011000011001",
   "011000011000",
   "011000011000",
   "011000010111",
   "011000010111",
   "011000010110",
   "011000010101",
   "011000010101",
   "011000010100",
   "011000010100",
   "011000010011",
   "011000010011",
   "011000010010",
   "011000010001",
   "011000010001",
   "011000010000",
   "011000010000",
   "011000001111",
   "011000001111",
   "011000001110",
   "011000001101",
   "011000001101",
   "011000001100",
   "011000001100",
   "011000001011",
   "011000001011",
   "011000001010",
   "011000001001",
   "011000001001",
   "011000001000",
   "011000001000",
   "011000000111",
   "011000000111",
   "011000000110",
   "011000000101",
   "011000000101",
   "011000000100",
   "011000000100",
   "011000000011",
   "011000000011",
   "011000000010",
   "011000000001",
   "011000000001",
   "011000000000",
   "011000000000",
   "010111111111",
   "010111111111",
   "010111111110",
   "010111111110",
   "010111111101",
   "010111111100",
   "010111111100",
   "010111111011",
   "010111111011",
   "010111111010",
   "010111111010",
   "010111111001",
   "010111111000",
   "010111111000",
   "010111110111",
   "010111110111",
   "010111110110",
   "010111110110",
   "010111110101",
   "010111110101",
   "010111110100",
   "010111110011",
   "010111110011",
   "010111110010",
   "010111110010",
   "010111110001",
   "010111110001",
   "010111110000",
   "010111110000",
   "010111101111",
   "010111101111",
   "010111101110",
   "010111101101",
   "010111101101",
   "010111101100",
   "010111101100",
   "010111101011",
   "010111101011",
   "010111101010",
   "010111101010",
   "010111101001",
   "010111101001",
   "010111101000",
   "010111100111",
   "010111100111",
   "010111100110",
   "010111100110",
   "010111100101",
   "010111100101",
   "010111100100",
   "010111100100",
   "010111100011",
   "010111100011",
   "010111100010",
   "010111100001",
   "010111100001",
   "010111100000",
   "010111100000",
   "010111011111",
   "010111011111",
   "010111011110",
   "010111011110",
   "010111011101",
   "010111011101",
   "010111011100",
   "010111011100",
   "010111011011",
   "010111011010",
   "010111011010",
   "010111011001",
   "010111011001",
   "010111011000",
   "010111011000",
   "010111010111",
   "010111010111",
   "010111010110",
   "010111010110",
   "010111010101",
   "010111010101",
   "010111010100",
   "010111010100",
   "010111010011",
   "010111010010",
   "010111010010",
   "010111010001",
   "010111010001",
   "010111010000",
   "010111010000",
   "010111001111",
   "010111001111",
   "010111001110",
   "010111001110",
   "010111001101",
   "010111001101",
   "010111001100",
   "010111001100",
   "010111001011",
   "010111001011",
   "010111001010",
   "010111001010",
   "010111001001",
   "010111001000",
   "010111001000",
   "010111000111",
   "010111000111",
   "010111000110",
   "010111000110",
   "010111000101",
   "010111000101",
   "010111000100",
   "010111000100",
   "010111000011",
   "010111000011",
   "010111000010",
   "010111000010",
   "010111000001",
   "010111000001",
   "010111000000",
   "010111000000",
   "010110111111",
   "010110111111",
   "010110111110",
   "010110111110",
   "010110111101",
   "010110111101",
   "010110111100",
   "010110111100",
   "010110111011",
   "010110111011",
   "010110111010",
   "010110111010",
   "010110111001",
   "010110111000",
   "010110111000",
   "010110110111",
   "010110110111",
   "010110110110",
   "010110110110",
   "010110110101",
   "010110110101",
   "010110110100",
   "010110110100",
   "010110110011",
   "010110110011",
   "010110110010",
   "010110110010",
   "010110110001",
   "010110110001",
   "010110110000",
   "010110110000",
   "010110101111",
   "010110101111",
   "010110101110",
   "010110101110",
   "010110101101",
   "010110101101",
   "010110101100",
   "010110101100",
   "010110101011",
   "010110101011",
   "010110101010",
   "010110101010",
   "010110101001",
   "010110101001",
   "010110101000",
   "010110101000",
   "010110100111",
   "010110100111",
   "010110100110",
   "010110100110",
   "010110100101",
   "010110100101",
   "010110100100",
   "010110100100",
   "010110100011",
   "010110100011",
   "010110100010",
   "010110100010",
   "010110100001",
   "010110100001",
   "010110100000",
   "010110100000",
   "010110011111",
   "010110011111",
   "010110011110",
   "010110011110",
   "010110011101",
   "010110011101",
   "010110011100",
   "010110011100",
   "010110011011",
   "010110011011",
   "010110011010",
   "010110011010",
   "010110011001",
   "010110011001",
   "010110011000",
   "010110011000",
   "010110011000",
   "010110010111",
   "010110010111",
   "010110010110",
   "010110010110",
   "010110010101",
   "010110010101",
   "010110010100",
   "010110010100",
   "010110010011",
   "010110010011",
   "010110010010",
   "010110010010",
   "010110010001",
   "010110010001",
   "010110010000",
   "010110010000",
   "010110001111",
   "010110001111",
   "010110001110",
   "010110001110",
   "010110001101",
   "010110001101",
   "010110001100",
   "010110001100",
   "010110001011",
   "010110001011",
   "010110001010",
   "010110001010",
   "010110001001",
   "010110001001",
   "010110001001",
   "010110001000",
   "010110001000",
   "010110000111",
   "010110000111",
   "010110000110",
   "010110000110",
   "010110000101",
   "010110000101",
   "010110000100",
   "010110000100",
   "010110000011",
   "010110000011",
   "010110000010",
   "010110000010",
   "010110000001",
   "010110000001",
   "010110000000",
   "010110000000",
   "010110000000",
   "010101111111",
   "010101111111",
   "010101111110",
   "010101111110",
   "010101111101",
   "010101111101",
   "010101111100",
   "010101111100",
   "010101111011",
   "010101111011",
   "010101111010",
   "010101111010",
   "010101111001",
   "010101111001",
   "010101111000",
   "010101111000",
   "010101111000",
   "010101110111",
   "010101110111",
   "010101110110",
   "010101110110",
   "010101110101",
   "010101110101",
   "010101110100",
   "010101110100",
   "010101110011",
   "010101110011",
   "010101110010",
   "010101110010",
   "010101110001",
   "010101110001",
   "010101110001",
   "010101110000",
   "010101110000",
   "010101101111",
   "010101101111",
   "010101101110",
   "010101101110",
   "010101101101",
   "010101101101",
   "010101101100",
   "010101101100",
   "010101101100",
   "010101101011",
   "010101101011",
   "010101101010",
   "010101101010",
   "010101101001",
   "010101101001",
   "010101101000",
   "010101101000",
   "010101100111",
   "010101100111",
   "010101100110",
   "010101100110",
   "010101100110",
   "010101100101",
   "010101100101",
   "010101100100",
   "010101100100",
   "010101100011",
   "010101100011",
   "010101100010",
   "010101100010",
   "010101100001",
   "010101100001",
   "010101100001",
   "010101100000",
   "010101100000",
   "010101011111",
   "010101011111",
   "010101011110",
   "010101011110",
   "010101011101",
   "010101011101",
   "010101011101",
   "010101011100",
   "010101011100",
   "010101011011",
   "010101011011",
   "010101011010",
   "010101011010",
   "010101011001",
   "010101011001",
   "010101011001",
   "010101011000",
   "010101011000",
   "010101010111",
   "010101010111",
   "010101010110",
   "101010101011",
   "101010101010",
   "101010101001",
   "101010101001",
   "101010101000",
   "101010100111",
   "101010100110",
   "101010100101",
   "101010100100",
   "101010100011",
   "101010100010",
   "101010100001",
   "101010100001",
   "101010100000",
   "101010011111",
   "101010011110",
   "101010011101",
   "101010011100",
   "101010011011",
   "101010011010",
   "101010011010",
   "101010011001",
   "101010011000",
   "101010010111",
   "101010010110",
   "101010010101",
   "101010010100",
   "101010010011",
   "101010010011",
   "101010010010",
   "101010010001",
   "101010010000",
   "101010001111",
   "101010001110",
   "101010001101",
   "101010001100",
   "101010001100",
   "101010001011",
   "101010001010",
   "101010001001",
   "101010001000",
   "101010000111",
   "101010000110",
   "101010000101",
   "101010000101",
   "101010000100",
   "101010000011",
   "101010000010",
   "101010000001",
   "101010000000",
   "101001111111",
   "101001111111",
   "101001111110",
   "101001111101",
   "101001111100",
   "101001111011",
   "101001111010",
   "101001111001",
   "101001111001",
   "101001111000",
   "101001110111",
   "101001110110",
   "101001110101",
   "101001110100",
   "101001110011",
   "101001110011",
   "101001110010",
   "101001110001",
   "101001110000",
   "101001101111",
   "101001101110",
   "101001101101",
   "101001101101",
   "101001101100",
   "101001101011",
   "101001101010",
   "101001101001",
   "101001101000",
   "101001101000",
   "101001100111",
   "101001100110",
   "101001100101",
   "101001100100",
   "101001100011",
   "101001100010",
   "101001100010",
   "101001100001",
   "101001100000",
   "101001011111",
   "101001011110",
   "101001011101",
   "101001011101",
   "101001011100",
   "101001011011",
   "101001011010",
   "101001011001",
   "101001011000",
   "101001011000",
   "101001010111",
   "101001010110",
   "101001010101",
   "101001010100",
   "101001010011",
   "101001010011",
   "101001010010",
   "101001010001",
   "101001010000",
   "101001001111",
   "101001001110",
   "101001001110",
   "101001001101",
   "101001001100",
   "101001001011",
   "101001001010",
   "101001001001",
   "101001001001",
   "101001001000",
   "101001000111",
   "101001000110",
   "101001000101",
   "101001000101",
   "101001000100",
   "101001000011",
   "101001000010",
   "101001000001",
   "101001000000",
   "101001000000",
   "101000111111",
   "101000111110",
   "101000111101",
   "101000111100",
   "101000111011",
   "101000111011",
   "101000111010",
   "101000111001",
   "101000111000",
   "101000110111",
   "101000110111",
   "101000110110",
   "101000110101",
   "101000110100",
   "101000110011",
   "101000110011",
   "101000110010",
   "101000110001",
   "101000110000",
   "101000101111",
   "101000101110",
   "101000101110",
   "101000101101",
   "101000101100",
   "101000101011",
   "101000101010",
   "101000101010",
   "101000101001",
   "101000101000",
   "101000100111",
   "101000100110",
   "101000100110",
   "101000100101",
   "101000100100",
   "101000100011",
   "101000100010",
   "101000100010",
   "101000100001",
   "101000100000",
   "101000011111",
   "101000011110",
   "101000011110",
   "101000011101",
   "101000011100",
   "101000011011",
   "101000011010",
   "101000011010",
   "101000011001",
   "101000011000",
   "101000010111",
   "101000010110",
   "101000010110",
   "101000010101",
   "101000010100",
   "101000010011",
   "101000010010",
   "101000010010",
   "101000010001",
   "101000010000",
   "101000001111",
   "101000001110",
   "101000001110",
   "101000001101",
   "101000001100",
   "101000001011",
   "101000001011",
   "101000001010",
   "101000001001",
   "101000001000",
   "101000000111",
   "101000000111",
   "101000000110",
   "101000000101",
   "101000000100",
   "101000000011",
   "101000000011",
   "101000000010",
   "101000000001",
   "101000000000",
   "101000000000",
   "100111111111",
   "100111111110",
   "100111111101",
   "100111111100",
   "100111111100",
   "100111111011",
   "100111111010",
   "100111111001",
   "100111111001",
   "100111111000",
   "100111110111",
   "100111110110",
   "100111110101",
   "100111110101",
   "100111110100",
   "100111110011",
   "100111110010",
   "100111110010",
   "100111110001",
   "100111110000",
   "100111101111",
   "100111101111",
   "100111101110",
   "100111101101",
   "100111101100",
   "100111101011",
   "100111101011",
   "100111101010",
   "100111101001",
   "100111101000",
   "100111101000",
   "100111100111",
   "100111100110",
   "100111100101",
   "100111100101",
   "100111100100",
   "100111100011",
   "100111100010",
   "100111100001",
   "100111100001",
   "100111100000",
   "100111011111",
   "100111011110",
   "100111011110",
   "100111011101",
   "100111011100",
   "100111011011",
   "100111011011",
   "100111011010",
   "100111011001",
   "100111011000",
   "100111011000",
   "100111010111",
   "100111010110",
   "100111010101",
   "100111010101",
   "100111010100",
   "100111010011",
   "100111010010",
   "100111010010",
   "100111010001",
   "100111010000",
   "100111001111",
   "100111001111",
   "100111001110",
   "100111001101",
   "100111001100",
   "100111001100",
   "100111001011",
   "100111001010",
   "100111001001",
   "100111001001",
   "100111001000",
   "100111000111",
   "100111000110",
   "100111000110",
   "100111000101",
   "100111000100",
   "100111000011",
   "100111000011",
   "100111000010",
   "100111000001",
   "100111000000",
   "100111000000",
   "100110111111",
   "100110111110",
   "100110111101",
   "100110111101",
   "100110111100",
   "100110111011",
   "100110111010",
   "100110111010",
   "100110111001",
   "100110111000",
   "100110110111",
   "100110110111",
   "100110110110",
   "100110110101",
   "100110110101",
   "100110110100",
   "100110110011",
   "100110110010",
   "100110110010",
   "100110110001",
   "100110110000",
   "100110101111",
   "100110101111",
   "100110101110",
   "100110101101",
   "100110101100",
   "100110101100",
   "100110101011",
   "100110101010",
   "100110101010",
   "100110101001",
   "100110101000",
   "100110100111",
   "100110100111",
   "100110100110",
   "100110100101",
   "100110100100",
   "100110100100",
   "100110100011",
   "100110100010",
   "100110100010",
   "100110100001",
   "100110100000",
   "100110011111",
   "100110011111",
   "100110011110",
   "100110011101",
   "100110011101",
   "100110011100",
   "100110011011",
   "100110011010",
   "100110011010",
   "100110011001",
   "100110011000",
   "100110010111",
   "100110010111",
   "100110010110",
   "100110010101",
   "100110010101",
   "100110010100",
   "100110010011",
   "100110010010",
   "100110010010",
   "100110010001",
   "100110010000",
   "100110010000",
   "100110001111",
   "100110001110",
   "100110001101",
   "100110001101",
   "100110001100",
   "100110001011",
   "100110001011",
   "100110001010",
   "100110001001",
   "100110001000",
   "100110001000",
   "100110000111",
   "100110000110",
   "100110000110",
   "100110000101",
   "100110000100",
   "100110000100",
   "100110000011",
   "100110000010",
   "100110000001",
   "100110000001",
   "100110000000",
   "100101111111",
   "100101111111",
   "100101111110",
   "100101111101",
   "100101111100",
   "100101111100",
   "100101111011",
   "100101111010",
   "100101111010",
   "100101111001",
   "100101111000",
   "100101111000",
   "100101110111",
   "100101110110",
   "100101110101",
   "100101110101",
   "100101110100",
   "100101110011",
   "100101110011",
   "100101110010",
   "100101110001",
   "100101110001",
   "100101110000",
   "100101101111",
   "100101101110",
   "100101101110",
   "100101101101",
   "100101101100",
   "100101101100",
   "100101101011",
   "100101101010",
   "100101101010",
   "100101101001",
   "100101101000",
   "100101101000",
   "100101100111",
   "100101100110",
   "100101100101",
   "100101100101",
   "100101100100",
   "100101100011",
   "100101100011",
   "100101100010",
   "100101100001",
   "100101100001",
   "100101100000",
   "100101011111",
   "100101011111",
   "100101011110",
   "100101011101",
   "100101011101",
   "100101011100",
   "100101011011",
   "100101011011",
   "100101011010",
   "100101011001",
   "100101011000",
   "100101011000",
   "100101010111",
   "100101010110",
   "100101010110",
   "100101010101",
   "100101010100",
   "100101010100",
   "100101010011",
   "100101010010",
   "100101010010",
   "100101010001",
   "100101010000",
   "100101010000",
   "100101001111",
   "100101001110",
   "100101001110",
   "100101001101",
   "100101001100",
   "100101001100",
   "100101001011",
   "100101001010",
   "100101001010",
   "100101001001",
   "100101001000",
   "100101001000",
   "100101000111",
   "100101000110",
   "100101000110",
   "100101000101",
   "100101000100",
   "100101000100",
   "100101000011",
   "100101000010",
   "100101000001",
   "100101000001",
   "100101000000",
   "100100111111",
   "100100111111",
   "100100111110",
   "100100111101",
   "100100111101",
   "100100111100",
   "100100111011",
   "100100111011",
   "100100111010",
   "100100111001",
   "100100111001",
   "100100111000",
   "100100111000",
   "100100110111",
   "100100110110",
   "100100110110",
   "100100110101",
   "100100110100",
   "100100110100",
   "100100110011",
   "100100110010",
   "100100110010",
   "100100110001",
   "100100110000",
   "100100110000",
   "100100101111",
   "100100101110",
   "100100101110",
   "100100101101",
   "100100101100",
   "100100101100",
   "100100101011",
   "100100101010",
   "100100101010",
   "100100101001",
   "100100101000",
   "100100101000",
   "100100100111",
   "100100100110",
   "100100100110",
   "100100100101",
   "100100100100",
   "100100100100",
   "100100100011",
   "100100100010",
   "100100100010",
   "100100100001",
   "100100100001",
   "100100100000",
   "100100011111",
   "100100011111",
   "100100011110",
   "100100011101",
   "100100011101",
   "100100011100",
   "100100011011",
   "100100011011",
   "100100011010",
   "100100011001",
   "100100011001",
   "100100011000",
   "100100010111",
   "100100010111",
   "100100010110",
   "100100010110",
   "100100010101",
   "100100010100",
   "100100010100",
   "100100010011",
   "100100010010",
   "100100010010",
   "100100010001",
   "100100010000",
   "100100010000",
   "100100001111",
   "100100001110",
   "100100001110",
   "100100001101",
   "100100001101",
   "100100001100",
   "100100001011",
   "100100001011",
   "100100001010",
   "100100001001",
   "100100001001",
   "100100001000",
   "100100000111",
   "100100000111",
   "100100000110",
   "100100000110",
   "100100000101",
   "100100000100",
   "100100000100",
   "100100000011",
   "100100000010",
   "100100000010",
   "100100000001",
   "100100000000",
   "100100000000",
   "100011111111",
   "100011111111",
   "100011111110",
   "100011111101",
   "100011111101",
   "100011111100",
   "100011111011",
   "100011111011",
   "100011111010",
   "100011111001",
   "100011111001",
   "100011111000",
   "100011111000",
   "100011110111",
   "100011110110",
   "100011110110",
   "100011110101",
   "100011110100",
   "100011110100",
   "100011110011",
   "100011110011",
   "100011110010",
   "100011110001",
   "100011110001",
   "100011110000",
   "100011101111",
   "100011101111",
   "100011101110",
   "100011101110",
   "100011101101",
   "100011101100",
   "100011101100",
   "100011101011",
   "100011101010",
   "100011101010",
   "100011101001",
   "100011101001",
   "100011101000",
   "100011100111",
   "100011100111",
   "100011100110",
   "100011100110",
   "100011100101",
   "100011100100",
   "100011100100",
   "100011100011",
   "100011100010",
   "100011100010",
   "100011100001",
   "100011100001",
   "100011100000",
   "100011011111",
   "100011011111",
   "100011011110",
   "100011011110",
   "100011011101",
   "100011011100",
   "100011011100",
   "100011011011",
   "100011011010",
   "100011011010",
   "100011011001",
   "100011011001",
   "100011011000",
   "100011010111",
   "100011010111",
   "100011010110",
   "100011010110",
   "100011010101",
   "100011010100",
   "100011010100",
   "100011010011",
   "100011010011",
   "100011010010",
   "100011010001",
   "100011010001",
   "100011010000",
   "100011010000",
   "100011001111",
   "100011001110",
   "100011001110",
   "100011001101",
   "100011001100",
   "100011001100",
   "100011001011",
   "100011001011",
   "100011001010",
   "100011001001",
   "100011001001",
   "100011001000",
   "100011001000",
   "100011000111",
   "100011000110",
   "100011000110",
   "100011000101",
   "100011000101",
   "100011000100",
   "100011000011",
   "100011000011",
   "100011000010",
   "100011000010",
   "100011000001",
   "100011000000",
   "100011000000",
   "100010111111",
   "100010111111",
   "100010111110",
   "100010111101",
   "100010111101",
   "100010111100",
   "100010111100",
   "100010111011",
   "100010111010",
   "100010111010",
   "100010111001",
   "100010111001",
   "100010111000",
   "100010111000",
   "100010110111",
   "100010110110",
   "100010110110",
   "100010110101",
   "100010110101",
   "100010110100",
   "100010110011",
   "100010110011",
   "100010110010",
   "100010110010",
   "100010110001",
   "100010110000",
   "100010110000",
   "100010101111",
   "100010101111",
   "100010101110",
   "100010101101",
   "100010101101",
   "100010101100",
   "100010101100",
   "100010101011",
   "100010101011",
   "100010101010",
   "100010101001",
   "100010101001",
   "100010101000",
   "100010101000",
   "100010100111",
   "100010100110",
   "100010100110",
   "100010100101",
   "100010100101",
   "100010100100",
   "100010100100",
   "100010100011",
   "100010100010",
   "100010100010",
   "100010100001",
   "100010100001",
   "100010100000",
   "100010011111",
   "100010011111",
   "100010011110",
   "100010011110",
   "100010011101",
   "100010011101",
   "100010011100",
   "100010011011",
   "100010011011",
   "100010011010",
   "100010011010",
   "100010011001",
   "100010011001",
   "100010011000",
   "100010010111",
   "100010010111",
   "100010010110",
   "100010010110",
   "100010010101",
   "100010010100",
   "100010010100",
   "100010010011",
   "100010010011",
   "100010010010",
   "100010010010",
   "100010010001",
   "100010010000",
   "100010010000",
   "100010001111",
   "100010001111",
   "100010001110",
   "100010001110",
   "100010001101",
   "100010001100",
   "100010001100",
   "100010001011",
   "100010001011",
   "100010001010",
   "100010001010",
   "100010001001",
   "100010001000",
   "100010001000",
   "100010000111",
   "100010000111",
   "100010000110",
   "100010000110",
   "100010000101",
   "100010000100",
   "100010000100",
   "100010000011",
   "100010000011",
   "100010000010",
   "100010000010",
   "100010000001",
   "100010000001",
   "100010000000",
   "100001111111",
   "100001111111",
   "100001111110",
   "100001111110",
   "100001111101",
   "100001111101",
   "100001111100",
   "100001111011",
   "100001111011",
   "100001111010",
   "100001111010",
   "100001111001",
   "100001111001",
   "100001111000",
   "100001111000",
   "100001110111",
   "100001110110",
   "100001110110",
   "100001110101",
   "100001110101",
   "100001110100",
   "100001110100",
   "100001110011",
   "100001110011",
   "100001110010",
   "100001110001",
   "100001110001",
   "100001110000",
   "100001110000",
   "100001101111",
   "100001101111",
   "100001101110",
   "100001101110",
   "100001101101",
   "100001101100",
   "100001101100",
   "100001101011",
   "100001101011",
   "100001101010",
   "100001101010",
   "100001101001",
   "100001101001",
   "100001101000",
   "100001100111",
   "100001100111",
   "100001100110",
   "100001100110",
   "100001100101",
   "100001100101",
   "100001100100",
   "100001100100",
   "100001100011",
   "100001100010",
   "100001100010",
   "100001100001",
   "100001100001",
   "100001100000",
   "100001100000",
   "100001011111",
   "100001011111",
   "100001011110",
   "100001011110",
   "100001011101",
   "100001011100",
   "100001011100",
   "100001011011",
   "100001011011",
   "100001011010",
   "100001011010",
   "100001011001",
   "100001011001",
   "100001011000",
   "100001011000",
   "100001010111",
   "100001010110",
   "100001010110",
   "100001010101",
   "100001010101",
   "100001010100",
   "100001010100",
   "100001010011",
   "100001010011",
   "100001010010",
   "100001010010",
   "100001010001",
   "100001010001",
   "100001010000",
   "100001001111",
   "100001001111",
   "100001001110",
   "100001001110",
   "100001001101",
   "100001001101",
   "100001001100",
   "100001001100",
   "100001001011",
   "100001001011",
   "100001001010",
   "100001001010",
   "100001001001",
   "100001001000",
   "100001001000",
   "100001000111",
   "100001000111",
   "100001000110",
   "100001000110",
   "100001000101",
   "100001000101",
   "100001000100",
   "100001000100",
   "100001000011",
   "100001000011",
   "100001000010",
   "100001000001",
   "100001000001",
   "100001000000",
   "100001000000",
   "100000111111",
   "100000111111",
   "100000111110",
   "100000111110",
   "100000111101",
   "100000111101",
   "100000111100",
   "100000111100",
   "100000111011",
   "100000111011",
   "100000111010",
   "100000111010",
   "100000111001",
   "100000111000",
   "100000111000",
   "100000110111",
   "100000110111",
   "100000110110",
   "100000110110",
   "100000110101",
   "100000110101",
   "100000110100",
   "100000110100",
   "100000110011",
   "100000110011",
   "100000110010",
   "100000110010",
   "100000110001",
   "100000110001",
   "100000110000",
   "100000110000",
   "100000101111",
   "100000101111",
   "100000101110",
   "100000101101",
   "100000101101",
   "100000101100",
   "100000101100",
   "100000101011",
   "100000101011",
   "100000101010",
   "100000101010",
   "100000101001",
   "100000101001",
   "100000101000",
   "100000101000",
   "100000100111",
   "100000100111",
   "100000100110",
   "100000100110",
   "100000100101",
   "100000100101",
   "100000100100",
   "100000100100",
   "100000100011",
   "100000100011",
   "100000100010",
   "100000100010",
   "100000100001",
   "100000100000",
   "100000100000",
   "100000011111",
   "100000011111",
   "100000011110",
   "100000011110",
   "100000011101",
   "100000011101",
   "100000011100",
   "100000011100",
   "100000011011",
   "100000011011",
   "100000011010",
   "100000011010",
   "100000011001",
   "100000011001",
   "100000011000",
   "100000011000",
   "100000010111",
   "100000010111",
   "100000010110",
   "100000010110",
   "100000010101",
   "100000010101",
   "100000010100",
   "100000010100",
   "100000010011",
   "100000010011",
   "100000010010",
   "100000010010",
   "100000010001",
   "100000010001",
   "100000010000",
   "100000010000",
   "100000001111",
   "100000001111",
   "100000001110",
   "100000001110",
   "100000001101",
   "100000001101",
   "100000001100",
   "100000001100",
   "100000001011",
   "100000001011",
   "100000001010",
   "100000001010",
   "100000001001",
   "100000001001",
   "100000001000",
   "100000001000",
   "100000000111",
   "100000000111",
   "100000000110",
   "100000000110",
   "100000000101",
   "100000000101",
   "100000000100",
   "100000000100",
   "100000000011",
   "100000000011",
   "100000000010",
   "100000000010",
   "100000000001",
      others => (others => '0'));
      	begin 
      return tmp;
      end init_rom;
	signal rom : memory_t := init_rom;
   signal Y0 :  std_logic_vector(11 downto 0);
begin
	process(clk)
   begin
   if(rising_edge(clk)) then
   	Y0 <= rom(  TO_INTEGER(unsigned(X))  );
   end if;
   end process;
    Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_67_f400_uid24
--                     (IntAdderClassical_67_f400_uid26)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_67_f400_uid24 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(66 downto 0);
          Y : in  std_logic_vector(66 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(66 downto 0)   );
end entity;

architecture arch of IntAdder_67_f400_uid24 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               IntMultiplier_UsingDSP_12_54_0_unsigned_uid11
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_12_54_0_unsigned_uid11 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          Y : in  std_logic_vector(53 downto 0);
          R : out  std_logic_vector(65 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_12_54_0_unsigned_uid11 is
   component IntAdder_67_f400_uid24 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(66 downto 0);
             Y : in  std_logic_vector(66 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(66 downto 0)   );
   end component;

signal XX_m12 :  std_logic_vector(53 downto 0);
signal YY_m12 :  std_logic_vector(11 downto 0);
signal DSP_bh13_ch0_0 :  std_logic_vector(40 downto 0);
signal heap_bh13_w65_0, heap_bh13_w65_0_d1 : std_logic;
signal heap_bh13_w64_0, heap_bh13_w64_0_d1 : std_logic;
signal heap_bh13_w63_0, heap_bh13_w63_0_d1 : std_logic;
signal heap_bh13_w62_0, heap_bh13_w62_0_d1 : std_logic;
signal heap_bh13_w61_0, heap_bh13_w61_0_d1 : std_logic;
signal heap_bh13_w60_0, heap_bh13_w60_0_d1 : std_logic;
signal heap_bh13_w59_0, heap_bh13_w59_0_d1 : std_logic;
signal heap_bh13_w58_0, heap_bh13_w58_0_d1 : std_logic;
signal heap_bh13_w57_0, heap_bh13_w57_0_d1 : std_logic;
signal heap_bh13_w56_0, heap_bh13_w56_0_d1 : std_logic;
signal heap_bh13_w55_0, heap_bh13_w55_0_d1 : std_logic;
signal heap_bh13_w54_0, heap_bh13_w54_0_d1 : std_logic;
signal heap_bh13_w53_0, heap_bh13_w53_0_d1 : std_logic;
signal heap_bh13_w52_0, heap_bh13_w52_0_d1 : std_logic;
signal heap_bh13_w51_0, heap_bh13_w51_0_d1 : std_logic;
signal heap_bh13_w50_0, heap_bh13_w50_0_d1 : std_logic;
signal heap_bh13_w49_0, heap_bh13_w49_0_d1 : std_logic;
signal heap_bh13_w48_0, heap_bh13_w48_0_d1 : std_logic;
signal heap_bh13_w47_0, heap_bh13_w47_0_d1 : std_logic;
signal heap_bh13_w46_0, heap_bh13_w46_0_d1 : std_logic;
signal heap_bh13_w45_0, heap_bh13_w45_0_d1 : std_logic;
signal heap_bh13_w44_0, heap_bh13_w44_0_d1 : std_logic;
signal heap_bh13_w43_0, heap_bh13_w43_0_d1 : std_logic;
signal heap_bh13_w42_0, heap_bh13_w42_0_d1 : std_logic;
signal heap_bh13_w41_0, heap_bh13_w41_0_d1 : std_logic;
signal heap_bh13_w40_0, heap_bh13_w40_0_d1 : std_logic;
signal heap_bh13_w39_0, heap_bh13_w39_0_d1 : std_logic;
signal heap_bh13_w38_0, heap_bh13_w38_0_d1 : std_logic;
signal heap_bh13_w37_0, heap_bh13_w37_0_d1 : std_logic;
signal heap_bh13_w36_0, heap_bh13_w36_0_d1 : std_logic;
signal heap_bh13_w35_0, heap_bh13_w35_0_d1 : std_logic;
signal heap_bh13_w34_0, heap_bh13_w34_0_d1 : std_logic;
signal heap_bh13_w33_0, heap_bh13_w33_0_d1 : std_logic;
signal heap_bh13_w32_0, heap_bh13_w32_0_d1 : std_logic;
signal heap_bh13_w31_0, heap_bh13_w31_0_d1 : std_logic;
signal heap_bh13_w30_0, heap_bh13_w30_0_d1 : std_logic;
signal heap_bh13_w29_0, heap_bh13_w29_0_d1 : std_logic;
signal heap_bh13_w28_0, heap_bh13_w28_0_d1 : std_logic;
signal heap_bh13_w27_0, heap_bh13_w27_0_d1 : std_logic;
signal heap_bh13_w26_0, heap_bh13_w26_0_d1 : std_logic;
signal heap_bh13_w25_0, heap_bh13_w25_0_d1 : std_logic;
signal DSP_bh13_ch1_0 :  std_logic_vector(40 downto 0);
signal heap_bh13_w41_1, heap_bh13_w41_1_d1 : std_logic;
signal heap_bh13_w40_1, heap_bh13_w40_1_d1 : std_logic;
signal heap_bh13_w39_1, heap_bh13_w39_1_d1 : std_logic;
signal heap_bh13_w38_1, heap_bh13_w38_1_d1 : std_logic;
signal heap_bh13_w37_1, heap_bh13_w37_1_d1 : std_logic;
signal heap_bh13_w36_1, heap_bh13_w36_1_d1 : std_logic;
signal heap_bh13_w35_1, heap_bh13_w35_1_d1 : std_logic;
signal heap_bh13_w34_1, heap_bh13_w34_1_d1 : std_logic;
signal heap_bh13_w33_1, heap_bh13_w33_1_d1 : std_logic;
signal heap_bh13_w32_1, heap_bh13_w32_1_d1 : std_logic;
signal heap_bh13_w31_1, heap_bh13_w31_1_d1 : std_logic;
signal heap_bh13_w30_1, heap_bh13_w30_1_d1 : std_logic;
signal heap_bh13_w29_1, heap_bh13_w29_1_d1 : std_logic;
signal heap_bh13_w28_1, heap_bh13_w28_1_d1 : std_logic;
signal heap_bh13_w27_1, heap_bh13_w27_1_d1 : std_logic;
signal heap_bh13_w26_1, heap_bh13_w26_1_d1 : std_logic;
signal heap_bh13_w25_1, heap_bh13_w25_1_d1 : std_logic;
signal heap_bh13_w24_0, heap_bh13_w24_0_d1 : std_logic;
signal heap_bh13_w23_0, heap_bh13_w23_0_d1 : std_logic;
signal heap_bh13_w22_0, heap_bh13_w22_0_d1 : std_logic;
signal heap_bh13_w21_0, heap_bh13_w21_0_d1 : std_logic;
signal heap_bh13_w20_0, heap_bh13_w20_0_d1 : std_logic;
signal heap_bh13_w19_0, heap_bh13_w19_0_d1 : std_logic;
signal heap_bh13_w18_0, heap_bh13_w18_0_d1 : std_logic;
signal heap_bh13_w17_0, heap_bh13_w17_0_d1 : std_logic;
signal heap_bh13_w16_0, heap_bh13_w16_0_d1 : std_logic;
signal heap_bh13_w15_0, heap_bh13_w15_0_d1 : std_logic;
signal heap_bh13_w14_0, heap_bh13_w14_0_d1 : std_logic;
signal heap_bh13_w13_0, heap_bh13_w13_0_d1 : std_logic;
signal heap_bh13_w12_0, heap_bh13_w12_0_d1 : std_logic;
signal heap_bh13_w11_0, heap_bh13_w11_0_d1 : std_logic;
signal heap_bh13_w10_0, heap_bh13_w10_0_d1 : std_logic;
signal heap_bh13_w9_0, heap_bh13_w9_0_d1 : std_logic;
signal heap_bh13_w8_0, heap_bh13_w8_0_d1 : std_logic;
signal heap_bh13_w7_0, heap_bh13_w7_0_d1 : std_logic;
signal heap_bh13_w6_0, heap_bh13_w6_0_d1 : std_logic;
signal heap_bh13_w5_0, heap_bh13_w5_0_d1 : std_logic;
signal heap_bh13_w4_0, heap_bh13_w4_0_d1 : std_logic;
signal heap_bh13_w3_0, heap_bh13_w3_0_d1 : std_logic;
signal heap_bh13_w2_0, heap_bh13_w2_0_d1 : std_logic;
signal heap_bh13_w1_0, heap_bh13_w1_0_d1 : std_logic;
signal DSP_bh13_ch2_0 :  std_logic_vector(40 downto 0);
signal heap_bh13_w17_1, heap_bh13_w17_1_d1 : std_logic;
signal heap_bh13_w16_1, heap_bh13_w16_1_d1 : std_logic;
signal heap_bh13_w15_1, heap_bh13_w15_1_d1 : std_logic;
signal heap_bh13_w14_1, heap_bh13_w14_1_d1 : std_logic;
signal heap_bh13_w13_1, heap_bh13_w13_1_d1 : std_logic;
signal heap_bh13_w12_1, heap_bh13_w12_1_d1 : std_logic;
signal heap_bh13_w11_1, heap_bh13_w11_1_d1 : std_logic;
signal heap_bh13_w10_1, heap_bh13_w10_1_d1 : std_logic;
signal heap_bh13_w9_1, heap_bh13_w9_1_d1 : std_logic;
signal heap_bh13_w8_1, heap_bh13_w8_1_d1 : std_logic;
signal heap_bh13_w7_1, heap_bh13_w7_1_d1 : std_logic;
signal heap_bh13_w6_1, heap_bh13_w6_1_d1 : std_logic;
signal heap_bh13_w5_1, heap_bh13_w5_1_d1 : std_logic;
signal heap_bh13_w4_1, heap_bh13_w4_1_d1 : std_logic;
signal heap_bh13_w3_1, heap_bh13_w3_1_d1 : std_logic;
signal heap_bh13_w2_1, heap_bh13_w2_1_d1 : std_logic;
signal heap_bh13_w1_1, heap_bh13_w1_1_d1 : std_logic;
signal heap_bh13_w0_0, heap_bh13_w0_0_d1 : std_logic;
signal finalAdderIn0_bh13 :  std_logic_vector(66 downto 0);
signal finalAdderIn1_bh13 :  std_logic_vector(66 downto 0);
signal finalAdderCin_bh13 : std_logic;
signal finalAdderOut_bh13 :  std_logic_vector(66 downto 0);
signal CompressionResult13 :  std_logic_vector(66 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            heap_bh13_w65_0_d1 <=  heap_bh13_w65_0;
            heap_bh13_w64_0_d1 <=  heap_bh13_w64_0;
            heap_bh13_w63_0_d1 <=  heap_bh13_w63_0;
            heap_bh13_w62_0_d1 <=  heap_bh13_w62_0;
            heap_bh13_w61_0_d1 <=  heap_bh13_w61_0;
            heap_bh13_w60_0_d1 <=  heap_bh13_w60_0;
            heap_bh13_w59_0_d1 <=  heap_bh13_w59_0;
            heap_bh13_w58_0_d1 <=  heap_bh13_w58_0;
            heap_bh13_w57_0_d1 <=  heap_bh13_w57_0;
            heap_bh13_w56_0_d1 <=  heap_bh13_w56_0;
            heap_bh13_w55_0_d1 <=  heap_bh13_w55_0;
            heap_bh13_w54_0_d1 <=  heap_bh13_w54_0;
            heap_bh13_w53_0_d1 <=  heap_bh13_w53_0;
            heap_bh13_w52_0_d1 <=  heap_bh13_w52_0;
            heap_bh13_w51_0_d1 <=  heap_bh13_w51_0;
            heap_bh13_w50_0_d1 <=  heap_bh13_w50_0;
            heap_bh13_w49_0_d1 <=  heap_bh13_w49_0;
            heap_bh13_w48_0_d1 <=  heap_bh13_w48_0;
            heap_bh13_w47_0_d1 <=  heap_bh13_w47_0;
            heap_bh13_w46_0_d1 <=  heap_bh13_w46_0;
            heap_bh13_w45_0_d1 <=  heap_bh13_w45_0;
            heap_bh13_w44_0_d1 <=  heap_bh13_w44_0;
            heap_bh13_w43_0_d1 <=  heap_bh13_w43_0;
            heap_bh13_w42_0_d1 <=  heap_bh13_w42_0;
            heap_bh13_w41_0_d1 <=  heap_bh13_w41_0;
            heap_bh13_w40_0_d1 <=  heap_bh13_w40_0;
            heap_bh13_w39_0_d1 <=  heap_bh13_w39_0;
            heap_bh13_w38_0_d1 <=  heap_bh13_w38_0;
            heap_bh13_w37_0_d1 <=  heap_bh13_w37_0;
            heap_bh13_w36_0_d1 <=  heap_bh13_w36_0;
            heap_bh13_w35_0_d1 <=  heap_bh13_w35_0;
            heap_bh13_w34_0_d1 <=  heap_bh13_w34_0;
            heap_bh13_w33_0_d1 <=  heap_bh13_w33_0;
            heap_bh13_w32_0_d1 <=  heap_bh13_w32_0;
            heap_bh13_w31_0_d1 <=  heap_bh13_w31_0;
            heap_bh13_w30_0_d1 <=  heap_bh13_w30_0;
            heap_bh13_w29_0_d1 <=  heap_bh13_w29_0;
            heap_bh13_w28_0_d1 <=  heap_bh13_w28_0;
            heap_bh13_w27_0_d1 <=  heap_bh13_w27_0;
            heap_bh13_w26_0_d1 <=  heap_bh13_w26_0;
            heap_bh13_w25_0_d1 <=  heap_bh13_w25_0;
            heap_bh13_w41_1_d1 <=  heap_bh13_w41_1;
            heap_bh13_w40_1_d1 <=  heap_bh13_w40_1;
            heap_bh13_w39_1_d1 <=  heap_bh13_w39_1;
            heap_bh13_w38_1_d1 <=  heap_bh13_w38_1;
            heap_bh13_w37_1_d1 <=  heap_bh13_w37_1;
            heap_bh13_w36_1_d1 <=  heap_bh13_w36_1;
            heap_bh13_w35_1_d1 <=  heap_bh13_w35_1;
            heap_bh13_w34_1_d1 <=  heap_bh13_w34_1;
            heap_bh13_w33_1_d1 <=  heap_bh13_w33_1;
            heap_bh13_w32_1_d1 <=  heap_bh13_w32_1;
            heap_bh13_w31_1_d1 <=  heap_bh13_w31_1;
            heap_bh13_w30_1_d1 <=  heap_bh13_w30_1;
            heap_bh13_w29_1_d1 <=  heap_bh13_w29_1;
            heap_bh13_w28_1_d1 <=  heap_bh13_w28_1;
            heap_bh13_w27_1_d1 <=  heap_bh13_w27_1;
            heap_bh13_w26_1_d1 <=  heap_bh13_w26_1;
            heap_bh13_w25_1_d1 <=  heap_bh13_w25_1;
            heap_bh13_w24_0_d1 <=  heap_bh13_w24_0;
            heap_bh13_w23_0_d1 <=  heap_bh13_w23_0;
            heap_bh13_w22_0_d1 <=  heap_bh13_w22_0;
            heap_bh13_w21_0_d1 <=  heap_bh13_w21_0;
            heap_bh13_w20_0_d1 <=  heap_bh13_w20_0;
            heap_bh13_w19_0_d1 <=  heap_bh13_w19_0;
            heap_bh13_w18_0_d1 <=  heap_bh13_w18_0;
            heap_bh13_w17_0_d1 <=  heap_bh13_w17_0;
            heap_bh13_w16_0_d1 <=  heap_bh13_w16_0;
            heap_bh13_w15_0_d1 <=  heap_bh13_w15_0;
            heap_bh13_w14_0_d1 <=  heap_bh13_w14_0;
            heap_bh13_w13_0_d1 <=  heap_bh13_w13_0;
            heap_bh13_w12_0_d1 <=  heap_bh13_w12_0;
            heap_bh13_w11_0_d1 <=  heap_bh13_w11_0;
            heap_bh13_w10_0_d1 <=  heap_bh13_w10_0;
            heap_bh13_w9_0_d1 <=  heap_bh13_w9_0;
            heap_bh13_w8_0_d1 <=  heap_bh13_w8_0;
            heap_bh13_w7_0_d1 <=  heap_bh13_w7_0;
            heap_bh13_w6_0_d1 <=  heap_bh13_w6_0;
            heap_bh13_w5_0_d1 <=  heap_bh13_w5_0;
            heap_bh13_w4_0_d1 <=  heap_bh13_w4_0;
            heap_bh13_w3_0_d1 <=  heap_bh13_w3_0;
            heap_bh13_w2_0_d1 <=  heap_bh13_w2_0;
            heap_bh13_w1_0_d1 <=  heap_bh13_w1_0;
            heap_bh13_w17_1_d1 <=  heap_bh13_w17_1;
            heap_bh13_w16_1_d1 <=  heap_bh13_w16_1;
            heap_bh13_w15_1_d1 <=  heap_bh13_w15_1;
            heap_bh13_w14_1_d1 <=  heap_bh13_w14_1;
            heap_bh13_w13_1_d1 <=  heap_bh13_w13_1;
            heap_bh13_w12_1_d1 <=  heap_bh13_w12_1;
            heap_bh13_w11_1_d1 <=  heap_bh13_w11_1;
            heap_bh13_w10_1_d1 <=  heap_bh13_w10_1;
            heap_bh13_w9_1_d1 <=  heap_bh13_w9_1;
            heap_bh13_w8_1_d1 <=  heap_bh13_w8_1;
            heap_bh13_w7_1_d1 <=  heap_bh13_w7_1;
            heap_bh13_w6_1_d1 <=  heap_bh13_w6_1;
            heap_bh13_w5_1_d1 <=  heap_bh13_w5_1;
            heap_bh13_w4_1_d1 <=  heap_bh13_w4_1;
            heap_bh13_w3_1_d1 <=  heap_bh13_w3_1;
            heap_bh13_w2_1_d1 <=  heap_bh13_w2_1;
            heap_bh13_w1_1_d1 <=  heap_bh13_w1_1;
            heap_bh13_w0_0_d1 <=  heap_bh13_w0_0;
         end if;
      end process;
   XX_m12 <= Y ;
   YY_m12 <= X ;
   
   -- Beginning of code generated by BitHeap::generateCompressorVHDL
   -- code generated by BitHeap::generateSupertileVHDL()
   ----------------Synchro barrier, entering cycle 0----------------
   DSP_bh13_ch0_0 <= ("" & XX_m12(53 downto 30) & "") * ("" & YY_m12(11 downto 0) & "00000");
   heap_bh13_w65_0 <= DSP_bh13_ch0_0(40); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w64_0 <= DSP_bh13_ch0_0(39); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w63_0 <= DSP_bh13_ch0_0(38); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w62_0 <= DSP_bh13_ch0_0(37); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w61_0 <= DSP_bh13_ch0_0(36); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w60_0 <= DSP_bh13_ch0_0(35); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w59_0 <= DSP_bh13_ch0_0(34); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w58_0 <= DSP_bh13_ch0_0(33); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w57_0 <= DSP_bh13_ch0_0(32); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w56_0 <= DSP_bh13_ch0_0(31); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w55_0 <= DSP_bh13_ch0_0(30); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w54_0 <= DSP_bh13_ch0_0(29); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w53_0 <= DSP_bh13_ch0_0(28); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w52_0 <= DSP_bh13_ch0_0(27); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w51_0 <= DSP_bh13_ch0_0(26); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w50_0 <= DSP_bh13_ch0_0(25); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w49_0 <= DSP_bh13_ch0_0(24); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w48_0 <= DSP_bh13_ch0_0(23); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w47_0 <= DSP_bh13_ch0_0(22); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w46_0 <= DSP_bh13_ch0_0(21); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w45_0 <= DSP_bh13_ch0_0(20); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w44_0 <= DSP_bh13_ch0_0(19); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w43_0 <= DSP_bh13_ch0_0(18); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w42_0 <= DSP_bh13_ch0_0(17); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w41_0 <= DSP_bh13_ch0_0(16); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w40_0 <= DSP_bh13_ch0_0(15); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w39_0 <= DSP_bh13_ch0_0(14); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w38_0 <= DSP_bh13_ch0_0(13); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w37_0 <= DSP_bh13_ch0_0(12); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w36_0 <= DSP_bh13_ch0_0(11); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w35_0 <= DSP_bh13_ch0_0(10); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w34_0 <= DSP_bh13_ch0_0(9); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w33_0 <= DSP_bh13_ch0_0(8); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w32_0 <= DSP_bh13_ch0_0(7); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w31_0 <= DSP_bh13_ch0_0(6); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w30_0 <= DSP_bh13_ch0_0(5); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w29_0 <= DSP_bh13_ch0_0(4); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w28_0 <= DSP_bh13_ch0_0(3); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w27_0 <= DSP_bh13_ch0_0(2); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w26_0 <= DSP_bh13_ch0_0(1); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w25_0 <= DSP_bh13_ch0_0(0); -- cycle= 0 cp= 1.638e-09
   ----------------Synchro barrier, entering cycle 0----------------
   DSP_bh13_ch1_0 <= ("" & XX_m12(29 downto 6) & "") * ("" & YY_m12(11 downto 0) & "00000");
   heap_bh13_w41_1 <= DSP_bh13_ch1_0(40); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w40_1 <= DSP_bh13_ch1_0(39); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w39_1 <= DSP_bh13_ch1_0(38); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w38_1 <= DSP_bh13_ch1_0(37); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w37_1 <= DSP_bh13_ch1_0(36); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w36_1 <= DSP_bh13_ch1_0(35); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w35_1 <= DSP_bh13_ch1_0(34); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w34_1 <= DSP_bh13_ch1_0(33); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w33_1 <= DSP_bh13_ch1_0(32); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w32_1 <= DSP_bh13_ch1_0(31); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w31_1 <= DSP_bh13_ch1_0(30); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w30_1 <= DSP_bh13_ch1_0(29); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w29_1 <= DSP_bh13_ch1_0(28); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w28_1 <= DSP_bh13_ch1_0(27); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w27_1 <= DSP_bh13_ch1_0(26); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w26_1 <= DSP_bh13_ch1_0(25); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w25_1 <= DSP_bh13_ch1_0(24); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w24_0 <= DSP_bh13_ch1_0(23); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w23_0 <= DSP_bh13_ch1_0(22); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w22_0 <= DSP_bh13_ch1_0(21); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w21_0 <= DSP_bh13_ch1_0(20); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w20_0 <= DSP_bh13_ch1_0(19); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w19_0 <= DSP_bh13_ch1_0(18); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w18_0 <= DSP_bh13_ch1_0(17); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w17_0 <= DSP_bh13_ch1_0(16); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w16_0 <= DSP_bh13_ch1_0(15); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w15_0 <= DSP_bh13_ch1_0(14); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w14_0 <= DSP_bh13_ch1_0(13); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w13_0 <= DSP_bh13_ch1_0(12); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w12_0 <= DSP_bh13_ch1_0(11); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w11_0 <= DSP_bh13_ch1_0(10); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w10_0 <= DSP_bh13_ch1_0(9); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w9_0 <= DSP_bh13_ch1_0(8); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w8_0 <= DSP_bh13_ch1_0(7); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w7_0 <= DSP_bh13_ch1_0(6); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w6_0 <= DSP_bh13_ch1_0(5); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w5_0 <= DSP_bh13_ch1_0(4); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w4_0 <= DSP_bh13_ch1_0(3); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w3_0 <= DSP_bh13_ch1_0(2); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w2_0 <= DSP_bh13_ch1_0(1); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w1_0 <= DSP_bh13_ch1_0(0); -- cycle= 0 cp= 1.638e-09
   ----------------Synchro barrier, entering cycle 0----------------
   DSP_bh13_ch2_0 <= ("" & XX_m12(5 downto 0) & "000000000000000000") * ("" & YY_m12(11 downto 0) & "00000");
   heap_bh13_w17_1 <= DSP_bh13_ch2_0(40); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w16_1 <= DSP_bh13_ch2_0(39); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w15_1 <= DSP_bh13_ch2_0(38); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w14_1 <= DSP_bh13_ch2_0(37); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w13_1 <= DSP_bh13_ch2_0(36); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w12_1 <= DSP_bh13_ch2_0(35); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w11_1 <= DSP_bh13_ch2_0(34); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w10_1 <= DSP_bh13_ch2_0(33); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w9_1 <= DSP_bh13_ch2_0(32); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w8_1 <= DSP_bh13_ch2_0(31); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w7_1 <= DSP_bh13_ch2_0(30); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w6_1 <= DSP_bh13_ch2_0(29); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w5_1 <= DSP_bh13_ch2_0(28); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w4_1 <= DSP_bh13_ch2_0(27); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w3_1 <= DSP_bh13_ch2_0(26); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w2_1 <= DSP_bh13_ch2_0(25); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w1_1 <= DSP_bh13_ch2_0(24); -- cycle= 0 cp= 1.638e-09
   heap_bh13_w0_0 <= DSP_bh13_ch2_0(23); -- cycle= 0 cp= 1.638e-09
   ----------------Synchro barrier, entering cycle 0----------------

   -- Adding the constant bits
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   finalAdderIn0_bh13 <= "0" & heap_bh13_w65_0_d1 & heap_bh13_w64_0_d1 & heap_bh13_w63_0_d1 & heap_bh13_w62_0_d1 & heap_bh13_w61_0_d1 & heap_bh13_w60_0_d1 & heap_bh13_w59_0_d1 & heap_bh13_w58_0_d1 & heap_bh13_w57_0_d1 & heap_bh13_w56_0_d1 & heap_bh13_w55_0_d1 & heap_bh13_w54_0_d1 & heap_bh13_w53_0_d1 & heap_bh13_w52_0_d1 & heap_bh13_w51_0_d1 & heap_bh13_w50_0_d1 & heap_bh13_w49_0_d1 & heap_bh13_w48_0_d1 & heap_bh13_w47_0_d1 & heap_bh13_w46_0_d1 & heap_bh13_w45_0_d1 & heap_bh13_w44_0_d1 & heap_bh13_w43_0_d1 & heap_bh13_w42_0_d1 & heap_bh13_w41_1_d1 & heap_bh13_w40_1_d1 & heap_bh13_w39_1_d1 & heap_bh13_w38_1_d1 & heap_bh13_w37_1_d1 & heap_bh13_w36_1_d1 & heap_bh13_w35_1_d1 & heap_bh13_w34_1_d1 & heap_bh13_w33_1_d1 & heap_bh13_w32_1_d1 & heap_bh13_w31_1_d1 & heap_bh13_w30_1_d1 & heap_bh13_w29_1_d1 & heap_bh13_w28_1_d1 & heap_bh13_w27_1_d1 & heap_bh13_w26_1_d1 & heap_bh13_w25_1_d1 & heap_bh13_w24_0_d1 & heap_bh13_w23_0_d1 & heap_bh13_w22_0_d1 & heap_bh13_w21_0_d1 & heap_bh13_w20_0_d1 & heap_bh13_w19_0_d1 & heap_bh13_w18_0_d1 & heap_bh13_w17_1_d1 & heap_bh13_w16_1_d1 & heap_bh13_w15_1_d1 & heap_bh13_w14_1_d1 & heap_bh13_w13_1_d1 & heap_bh13_w12_1_d1 & heap_bh13_w11_1_d1 & heap_bh13_w10_1_d1 & heap_bh13_w9_1_d1 & heap_bh13_w8_1_d1 & heap_bh13_w7_1_d1 & heap_bh13_w6_1_d1 & heap_bh13_w5_1_d1 & heap_bh13_w4_1_d1 & heap_bh13_w3_1_d1 & heap_bh13_w2_1_d1 & heap_bh13_w1_1_d1 & heap_bh13_w0_0_d1;
   finalAdderIn1_bh13 <= "0" & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh13_w41_0_d1 & heap_bh13_w40_0_d1 & heap_bh13_w39_0_d1 & heap_bh13_w38_0_d1 & heap_bh13_w37_0_d1 & heap_bh13_w36_0_d1 & heap_bh13_w35_0_d1 & heap_bh13_w34_0_d1 & heap_bh13_w33_0_d1 & heap_bh13_w32_0_d1 & heap_bh13_w31_0_d1 & heap_bh13_w30_0_d1 & heap_bh13_w29_0_d1 & heap_bh13_w28_0_d1 & heap_bh13_w27_0_d1 & heap_bh13_w26_0_d1 & heap_bh13_w25_0_d1 & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh13_w17_0_d1 & heap_bh13_w16_0_d1 & heap_bh13_w15_0_d1 & heap_bh13_w14_0_d1 & heap_bh13_w13_0_d1 & heap_bh13_w12_0_d1 & heap_bh13_w11_0_d1 & heap_bh13_w10_0_d1 & heap_bh13_w9_0_d1 & heap_bh13_w8_0_d1 & heap_bh13_w7_0_d1 & heap_bh13_w6_0_d1 & heap_bh13_w5_0_d1 & heap_bh13_w4_0_d1 & heap_bh13_w3_0_d1 & heap_bh13_w2_0_d1 & heap_bh13_w1_0_d1 & '0';
   finalAdderCin_bh13 <= '0';
   Adder_final13_0: IntAdder_67_f400_uid24  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => finalAdderCin_bh13,
                 R => finalAdderOut_bh13   ,
                 X => finalAdderIn0_bh13,
                 Y => finalAdderIn1_bh13);
   -- concatenate all the compressed chunks
   CompressionResult13 <= finalAdderOut_bh13;
   -- End of code generated by BitHeap::generateCompressorVHDL
   R <= CompressionResult13(65 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_65_f400_uid45
--                     (IntAdderClassical_65_f400_uid47)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_65_f400_uid45 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(64 downto 0);
          Y : in  std_logic_vector(64 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(64 downto 0)   );
end entity;

architecture arch of IntAdder_65_f400_uid45 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                IntMultiplier_UsingDSP_9_55_0_unsigned_uid32
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_9_55_0_unsigned_uid32 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(8 downto 0);
          Y : in  std_logic_vector(54 downto 0);
          R : out  std_logic_vector(63 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_9_55_0_unsigned_uid32 is
   component IntAdder_65_f400_uid45 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(64 downto 0);
             Y : in  std_logic_vector(64 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(64 downto 0)   );
   end component;

signal XX_m33 :  std_logic_vector(54 downto 0);
signal YY_m33 :  std_logic_vector(8 downto 0);
signal DSP_bh34_ch0_0 :  std_logic_vector(40 downto 0);
signal heap_bh34_w63_0, heap_bh34_w63_0_d1 : std_logic;
signal heap_bh34_w62_0, heap_bh34_w62_0_d1 : std_logic;
signal heap_bh34_w61_0, heap_bh34_w61_0_d1 : std_logic;
signal heap_bh34_w60_0, heap_bh34_w60_0_d1 : std_logic;
signal heap_bh34_w59_0, heap_bh34_w59_0_d1 : std_logic;
signal heap_bh34_w58_0, heap_bh34_w58_0_d1 : std_logic;
signal heap_bh34_w57_0, heap_bh34_w57_0_d1 : std_logic;
signal heap_bh34_w56_0, heap_bh34_w56_0_d1 : std_logic;
signal heap_bh34_w55_0, heap_bh34_w55_0_d1 : std_logic;
signal heap_bh34_w54_0, heap_bh34_w54_0_d1 : std_logic;
signal heap_bh34_w53_0, heap_bh34_w53_0_d1 : std_logic;
signal heap_bh34_w52_0, heap_bh34_w52_0_d1 : std_logic;
signal heap_bh34_w51_0, heap_bh34_w51_0_d1 : std_logic;
signal heap_bh34_w50_0, heap_bh34_w50_0_d1 : std_logic;
signal heap_bh34_w49_0, heap_bh34_w49_0_d1 : std_logic;
signal heap_bh34_w48_0, heap_bh34_w48_0_d1 : std_logic;
signal heap_bh34_w47_0, heap_bh34_w47_0_d1 : std_logic;
signal heap_bh34_w46_0, heap_bh34_w46_0_d1 : std_logic;
signal heap_bh34_w45_0, heap_bh34_w45_0_d1 : std_logic;
signal heap_bh34_w44_0, heap_bh34_w44_0_d1 : std_logic;
signal heap_bh34_w43_0, heap_bh34_w43_0_d1 : std_logic;
signal heap_bh34_w42_0, heap_bh34_w42_0_d1 : std_logic;
signal heap_bh34_w41_0, heap_bh34_w41_0_d1 : std_logic;
signal heap_bh34_w40_0, heap_bh34_w40_0_d1 : std_logic;
signal heap_bh34_w39_0, heap_bh34_w39_0_d1 : std_logic;
signal heap_bh34_w38_0, heap_bh34_w38_0_d1 : std_logic;
signal heap_bh34_w37_0, heap_bh34_w37_0_d1 : std_logic;
signal heap_bh34_w36_0, heap_bh34_w36_0_d1 : std_logic;
signal heap_bh34_w35_0, heap_bh34_w35_0_d1 : std_logic;
signal heap_bh34_w34_0, heap_bh34_w34_0_d1 : std_logic;
signal heap_bh34_w33_0, heap_bh34_w33_0_d1 : std_logic;
signal heap_bh34_w32_0, heap_bh34_w32_0_d1 : std_logic;
signal heap_bh34_w31_0, heap_bh34_w31_0_d1 : std_logic;
signal heap_bh34_w30_0, heap_bh34_w30_0_d1 : std_logic;
signal heap_bh34_w29_0, heap_bh34_w29_0_d1 : std_logic;
signal heap_bh34_w28_0, heap_bh34_w28_0_d1 : std_logic;
signal heap_bh34_w27_0, heap_bh34_w27_0_d1 : std_logic;
signal heap_bh34_w26_0, heap_bh34_w26_0_d1 : std_logic;
signal heap_bh34_w25_0, heap_bh34_w25_0_d1 : std_logic;
signal heap_bh34_w24_0, heap_bh34_w24_0_d1 : std_logic;
signal heap_bh34_w23_0, heap_bh34_w23_0_d1 : std_logic;
signal DSP_bh34_ch1_0 :  std_logic_vector(40 downto 0);
signal heap_bh34_w39_1, heap_bh34_w39_1_d1 : std_logic;
signal heap_bh34_w38_1, heap_bh34_w38_1_d1 : std_logic;
signal heap_bh34_w37_1, heap_bh34_w37_1_d1 : std_logic;
signal heap_bh34_w36_1, heap_bh34_w36_1_d1 : std_logic;
signal heap_bh34_w35_1, heap_bh34_w35_1_d1 : std_logic;
signal heap_bh34_w34_1, heap_bh34_w34_1_d1 : std_logic;
signal heap_bh34_w33_1, heap_bh34_w33_1_d1 : std_logic;
signal heap_bh34_w32_1, heap_bh34_w32_1_d1 : std_logic;
signal heap_bh34_w31_1, heap_bh34_w31_1_d1 : std_logic;
signal heap_bh34_w30_1, heap_bh34_w30_1_d1 : std_logic;
signal heap_bh34_w29_1, heap_bh34_w29_1_d1 : std_logic;
signal heap_bh34_w28_1, heap_bh34_w28_1_d1 : std_logic;
signal heap_bh34_w27_1, heap_bh34_w27_1_d1 : std_logic;
signal heap_bh34_w26_1, heap_bh34_w26_1_d1 : std_logic;
signal heap_bh34_w25_1, heap_bh34_w25_1_d1 : std_logic;
signal heap_bh34_w24_1, heap_bh34_w24_1_d1 : std_logic;
signal heap_bh34_w23_1, heap_bh34_w23_1_d1 : std_logic;
signal heap_bh34_w22_0, heap_bh34_w22_0_d1 : std_logic;
signal heap_bh34_w21_0, heap_bh34_w21_0_d1 : std_logic;
signal heap_bh34_w20_0, heap_bh34_w20_0_d1 : std_logic;
signal heap_bh34_w19_0, heap_bh34_w19_0_d1 : std_logic;
signal heap_bh34_w18_0, heap_bh34_w18_0_d1 : std_logic;
signal heap_bh34_w17_0, heap_bh34_w17_0_d1 : std_logic;
signal heap_bh34_w16_0, heap_bh34_w16_0_d1 : std_logic;
signal heap_bh34_w15_0, heap_bh34_w15_0_d1 : std_logic;
signal heap_bh34_w14_0, heap_bh34_w14_0_d1 : std_logic;
signal heap_bh34_w13_0, heap_bh34_w13_0_d1 : std_logic;
signal heap_bh34_w12_0, heap_bh34_w12_0_d1 : std_logic;
signal heap_bh34_w11_0, heap_bh34_w11_0_d1 : std_logic;
signal heap_bh34_w10_0, heap_bh34_w10_0_d1 : std_logic;
signal heap_bh34_w9_0, heap_bh34_w9_0_d1 : std_logic;
signal heap_bh34_w8_0, heap_bh34_w8_0_d1 : std_logic;
signal heap_bh34_w7_0, heap_bh34_w7_0_d1 : std_logic;
signal heap_bh34_w6_0, heap_bh34_w6_0_d1 : std_logic;
signal heap_bh34_w5_0, heap_bh34_w5_0_d1 : std_logic;
signal heap_bh34_w4_0, heap_bh34_w4_0_d1 : std_logic;
signal heap_bh34_w3_0, heap_bh34_w3_0_d1 : std_logic;
signal heap_bh34_w2_0, heap_bh34_w2_0_d1 : std_logic;
signal heap_bh34_w1_0, heap_bh34_w1_0_d1 : std_logic;
signal heap_bh34_w0_0, heap_bh34_w0_0_d1 : std_logic;
signal DSP_bh34_ch2_0 :  std_logic_vector(40 downto 0);
signal heap_bh34_w15_1, heap_bh34_w15_1_d1 : std_logic;
signal heap_bh34_w14_1, heap_bh34_w14_1_d1 : std_logic;
signal heap_bh34_w13_1, heap_bh34_w13_1_d1 : std_logic;
signal heap_bh34_w12_1, heap_bh34_w12_1_d1 : std_logic;
signal heap_bh34_w11_1, heap_bh34_w11_1_d1 : std_logic;
signal heap_bh34_w10_1, heap_bh34_w10_1_d1 : std_logic;
signal heap_bh34_w9_1, heap_bh34_w9_1_d1 : std_logic;
signal heap_bh34_w8_1, heap_bh34_w8_1_d1 : std_logic;
signal heap_bh34_w7_1, heap_bh34_w7_1_d1 : std_logic;
signal heap_bh34_w6_1, heap_bh34_w6_1_d1 : std_logic;
signal heap_bh34_w5_1, heap_bh34_w5_1_d1 : std_logic;
signal heap_bh34_w4_1, heap_bh34_w4_1_d1 : std_logic;
signal heap_bh34_w3_1, heap_bh34_w3_1_d1 : std_logic;
signal heap_bh34_w2_1, heap_bh34_w2_1_d1 : std_logic;
signal heap_bh34_w1_1, heap_bh34_w1_1_d1 : std_logic;
signal heap_bh34_w0_1, heap_bh34_w0_1_d1 : std_logic;
signal finalAdderIn0_bh34 :  std_logic_vector(64 downto 0);
signal finalAdderIn1_bh34 :  std_logic_vector(64 downto 0);
signal finalAdderCin_bh34 : std_logic;
signal finalAdderOut_bh34 :  std_logic_vector(64 downto 0);
signal CompressionResult34 :  std_logic_vector(64 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            heap_bh34_w63_0_d1 <=  heap_bh34_w63_0;
            heap_bh34_w62_0_d1 <=  heap_bh34_w62_0;
            heap_bh34_w61_0_d1 <=  heap_bh34_w61_0;
            heap_bh34_w60_0_d1 <=  heap_bh34_w60_0;
            heap_bh34_w59_0_d1 <=  heap_bh34_w59_0;
            heap_bh34_w58_0_d1 <=  heap_bh34_w58_0;
            heap_bh34_w57_0_d1 <=  heap_bh34_w57_0;
            heap_bh34_w56_0_d1 <=  heap_bh34_w56_0;
            heap_bh34_w55_0_d1 <=  heap_bh34_w55_0;
            heap_bh34_w54_0_d1 <=  heap_bh34_w54_0;
            heap_bh34_w53_0_d1 <=  heap_bh34_w53_0;
            heap_bh34_w52_0_d1 <=  heap_bh34_w52_0;
            heap_bh34_w51_0_d1 <=  heap_bh34_w51_0;
            heap_bh34_w50_0_d1 <=  heap_bh34_w50_0;
            heap_bh34_w49_0_d1 <=  heap_bh34_w49_0;
            heap_bh34_w48_0_d1 <=  heap_bh34_w48_0;
            heap_bh34_w47_0_d1 <=  heap_bh34_w47_0;
            heap_bh34_w46_0_d1 <=  heap_bh34_w46_0;
            heap_bh34_w45_0_d1 <=  heap_bh34_w45_0;
            heap_bh34_w44_0_d1 <=  heap_bh34_w44_0;
            heap_bh34_w43_0_d1 <=  heap_bh34_w43_0;
            heap_bh34_w42_0_d1 <=  heap_bh34_w42_0;
            heap_bh34_w41_0_d1 <=  heap_bh34_w41_0;
            heap_bh34_w40_0_d1 <=  heap_bh34_w40_0;
            heap_bh34_w39_0_d1 <=  heap_bh34_w39_0;
            heap_bh34_w38_0_d1 <=  heap_bh34_w38_0;
            heap_bh34_w37_0_d1 <=  heap_bh34_w37_0;
            heap_bh34_w36_0_d1 <=  heap_bh34_w36_0;
            heap_bh34_w35_0_d1 <=  heap_bh34_w35_0;
            heap_bh34_w34_0_d1 <=  heap_bh34_w34_0;
            heap_bh34_w33_0_d1 <=  heap_bh34_w33_0;
            heap_bh34_w32_0_d1 <=  heap_bh34_w32_0;
            heap_bh34_w31_0_d1 <=  heap_bh34_w31_0;
            heap_bh34_w30_0_d1 <=  heap_bh34_w30_0;
            heap_bh34_w29_0_d1 <=  heap_bh34_w29_0;
            heap_bh34_w28_0_d1 <=  heap_bh34_w28_0;
            heap_bh34_w27_0_d1 <=  heap_bh34_w27_0;
            heap_bh34_w26_0_d1 <=  heap_bh34_w26_0;
            heap_bh34_w25_0_d1 <=  heap_bh34_w25_0;
            heap_bh34_w24_0_d1 <=  heap_bh34_w24_0;
            heap_bh34_w23_0_d1 <=  heap_bh34_w23_0;
            heap_bh34_w39_1_d1 <=  heap_bh34_w39_1;
            heap_bh34_w38_1_d1 <=  heap_bh34_w38_1;
            heap_bh34_w37_1_d1 <=  heap_bh34_w37_1;
            heap_bh34_w36_1_d1 <=  heap_bh34_w36_1;
            heap_bh34_w35_1_d1 <=  heap_bh34_w35_1;
            heap_bh34_w34_1_d1 <=  heap_bh34_w34_1;
            heap_bh34_w33_1_d1 <=  heap_bh34_w33_1;
            heap_bh34_w32_1_d1 <=  heap_bh34_w32_1;
            heap_bh34_w31_1_d1 <=  heap_bh34_w31_1;
            heap_bh34_w30_1_d1 <=  heap_bh34_w30_1;
            heap_bh34_w29_1_d1 <=  heap_bh34_w29_1;
            heap_bh34_w28_1_d1 <=  heap_bh34_w28_1;
            heap_bh34_w27_1_d1 <=  heap_bh34_w27_1;
            heap_bh34_w26_1_d1 <=  heap_bh34_w26_1;
            heap_bh34_w25_1_d1 <=  heap_bh34_w25_1;
            heap_bh34_w24_1_d1 <=  heap_bh34_w24_1;
            heap_bh34_w23_1_d1 <=  heap_bh34_w23_1;
            heap_bh34_w22_0_d1 <=  heap_bh34_w22_0;
            heap_bh34_w21_0_d1 <=  heap_bh34_w21_0;
            heap_bh34_w20_0_d1 <=  heap_bh34_w20_0;
            heap_bh34_w19_0_d1 <=  heap_bh34_w19_0;
            heap_bh34_w18_0_d1 <=  heap_bh34_w18_0;
            heap_bh34_w17_0_d1 <=  heap_bh34_w17_0;
            heap_bh34_w16_0_d1 <=  heap_bh34_w16_0;
            heap_bh34_w15_0_d1 <=  heap_bh34_w15_0;
            heap_bh34_w14_0_d1 <=  heap_bh34_w14_0;
            heap_bh34_w13_0_d1 <=  heap_bh34_w13_0;
            heap_bh34_w12_0_d1 <=  heap_bh34_w12_0;
            heap_bh34_w11_0_d1 <=  heap_bh34_w11_0;
            heap_bh34_w10_0_d1 <=  heap_bh34_w10_0;
            heap_bh34_w9_0_d1 <=  heap_bh34_w9_0;
            heap_bh34_w8_0_d1 <=  heap_bh34_w8_0;
            heap_bh34_w7_0_d1 <=  heap_bh34_w7_0;
            heap_bh34_w6_0_d1 <=  heap_bh34_w6_0;
            heap_bh34_w5_0_d1 <=  heap_bh34_w5_0;
            heap_bh34_w4_0_d1 <=  heap_bh34_w4_0;
            heap_bh34_w3_0_d1 <=  heap_bh34_w3_0;
            heap_bh34_w2_0_d1 <=  heap_bh34_w2_0;
            heap_bh34_w1_0_d1 <=  heap_bh34_w1_0;
            heap_bh34_w0_0_d1 <=  heap_bh34_w0_0;
            heap_bh34_w15_1_d1 <=  heap_bh34_w15_1;
            heap_bh34_w14_1_d1 <=  heap_bh34_w14_1;
            heap_bh34_w13_1_d1 <=  heap_bh34_w13_1;
            heap_bh34_w12_1_d1 <=  heap_bh34_w12_1;
            heap_bh34_w11_1_d1 <=  heap_bh34_w11_1;
            heap_bh34_w10_1_d1 <=  heap_bh34_w10_1;
            heap_bh34_w9_1_d1 <=  heap_bh34_w9_1;
            heap_bh34_w8_1_d1 <=  heap_bh34_w8_1;
            heap_bh34_w7_1_d1 <=  heap_bh34_w7_1;
            heap_bh34_w6_1_d1 <=  heap_bh34_w6_1;
            heap_bh34_w5_1_d1 <=  heap_bh34_w5_1;
            heap_bh34_w4_1_d1 <=  heap_bh34_w4_1;
            heap_bh34_w3_1_d1 <=  heap_bh34_w3_1;
            heap_bh34_w2_1_d1 <=  heap_bh34_w2_1;
            heap_bh34_w1_1_d1 <=  heap_bh34_w1_1;
            heap_bh34_w0_1_d1 <=  heap_bh34_w0_1;
         end if;
      end process;
   XX_m33 <= Y ;
   YY_m33 <= X ;
   
   -- Beginning of code generated by BitHeap::generateCompressorVHDL
   -- code generated by BitHeap::generateSupertileVHDL()
   ----------------Synchro barrier, entering cycle 0----------------
   DSP_bh34_ch0_0 <= ("" & XX_m33(54 downto 31) & "") * ("" & YY_m33(8 downto 0) & "00000000");
   heap_bh34_w63_0 <= DSP_bh34_ch0_0(40); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w62_0 <= DSP_bh34_ch0_0(39); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w61_0 <= DSP_bh34_ch0_0(38); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w60_0 <= DSP_bh34_ch0_0(37); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w59_0 <= DSP_bh34_ch0_0(36); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w58_0 <= DSP_bh34_ch0_0(35); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w57_0 <= DSP_bh34_ch0_0(34); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w56_0 <= DSP_bh34_ch0_0(33); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w55_0 <= DSP_bh34_ch0_0(32); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w54_0 <= DSP_bh34_ch0_0(31); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w53_0 <= DSP_bh34_ch0_0(30); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w52_0 <= DSP_bh34_ch0_0(29); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w51_0 <= DSP_bh34_ch0_0(28); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w50_0 <= DSP_bh34_ch0_0(27); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w49_0 <= DSP_bh34_ch0_0(26); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w48_0 <= DSP_bh34_ch0_0(25); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w47_0 <= DSP_bh34_ch0_0(24); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w46_0 <= DSP_bh34_ch0_0(23); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w45_0 <= DSP_bh34_ch0_0(22); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w44_0 <= DSP_bh34_ch0_0(21); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w43_0 <= DSP_bh34_ch0_0(20); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w42_0 <= DSP_bh34_ch0_0(19); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w41_0 <= DSP_bh34_ch0_0(18); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w40_0 <= DSP_bh34_ch0_0(17); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w39_0 <= DSP_bh34_ch0_0(16); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w38_0 <= DSP_bh34_ch0_0(15); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w37_0 <= DSP_bh34_ch0_0(14); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w36_0 <= DSP_bh34_ch0_0(13); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w35_0 <= DSP_bh34_ch0_0(12); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w34_0 <= DSP_bh34_ch0_0(11); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w33_0 <= DSP_bh34_ch0_0(10); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w32_0 <= DSP_bh34_ch0_0(9); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w31_0 <= DSP_bh34_ch0_0(8); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w30_0 <= DSP_bh34_ch0_0(7); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w29_0 <= DSP_bh34_ch0_0(6); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w28_0 <= DSP_bh34_ch0_0(5); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w27_0 <= DSP_bh34_ch0_0(4); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w26_0 <= DSP_bh34_ch0_0(3); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w25_0 <= DSP_bh34_ch0_0(2); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w24_0 <= DSP_bh34_ch0_0(1); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w23_0 <= DSP_bh34_ch0_0(0); -- cycle= 0 cp= 1.638e-09
   ----------------Synchro barrier, entering cycle 0----------------
   DSP_bh34_ch1_0 <= ("" & XX_m33(30 downto 7) & "") * ("" & YY_m33(8 downto 0) & "00000000");
   heap_bh34_w39_1 <= DSP_bh34_ch1_0(40); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w38_1 <= DSP_bh34_ch1_0(39); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w37_1 <= DSP_bh34_ch1_0(38); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w36_1 <= DSP_bh34_ch1_0(37); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w35_1 <= DSP_bh34_ch1_0(36); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w34_1 <= DSP_bh34_ch1_0(35); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w33_1 <= DSP_bh34_ch1_0(34); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w32_1 <= DSP_bh34_ch1_0(33); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w31_1 <= DSP_bh34_ch1_0(32); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w30_1 <= DSP_bh34_ch1_0(31); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w29_1 <= DSP_bh34_ch1_0(30); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w28_1 <= DSP_bh34_ch1_0(29); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w27_1 <= DSP_bh34_ch1_0(28); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w26_1 <= DSP_bh34_ch1_0(27); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w25_1 <= DSP_bh34_ch1_0(26); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w24_1 <= DSP_bh34_ch1_0(25); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w23_1 <= DSP_bh34_ch1_0(24); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w22_0 <= DSP_bh34_ch1_0(23); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w21_0 <= DSP_bh34_ch1_0(22); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w20_0 <= DSP_bh34_ch1_0(21); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w19_0 <= DSP_bh34_ch1_0(20); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w18_0 <= DSP_bh34_ch1_0(19); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w17_0 <= DSP_bh34_ch1_0(18); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w16_0 <= DSP_bh34_ch1_0(17); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w15_0 <= DSP_bh34_ch1_0(16); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w14_0 <= DSP_bh34_ch1_0(15); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w13_0 <= DSP_bh34_ch1_0(14); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w12_0 <= DSP_bh34_ch1_0(13); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w11_0 <= DSP_bh34_ch1_0(12); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w10_0 <= DSP_bh34_ch1_0(11); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w9_0 <= DSP_bh34_ch1_0(10); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w8_0 <= DSP_bh34_ch1_0(9); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w7_0 <= DSP_bh34_ch1_0(8); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w6_0 <= DSP_bh34_ch1_0(7); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w5_0 <= DSP_bh34_ch1_0(6); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w4_0 <= DSP_bh34_ch1_0(5); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w3_0 <= DSP_bh34_ch1_0(4); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w2_0 <= DSP_bh34_ch1_0(3); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w1_0 <= DSP_bh34_ch1_0(2); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w0_0 <= DSP_bh34_ch1_0(1); -- cycle= 0 cp= 1.638e-09
   ----------------Synchro barrier, entering cycle 0----------------
   DSP_bh34_ch2_0 <= ("" & XX_m33(6 downto 0) & "00000000000000000") * ("" & YY_m33(8 downto 0) & "00000000");
   heap_bh34_w15_1 <= DSP_bh34_ch2_0(40); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w14_1 <= DSP_bh34_ch2_0(39); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w13_1 <= DSP_bh34_ch2_0(38); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w12_1 <= DSP_bh34_ch2_0(37); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w11_1 <= DSP_bh34_ch2_0(36); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w10_1 <= DSP_bh34_ch2_0(35); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w9_1 <= DSP_bh34_ch2_0(34); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w8_1 <= DSP_bh34_ch2_0(33); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w7_1 <= DSP_bh34_ch2_0(32); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w6_1 <= DSP_bh34_ch2_0(31); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w5_1 <= DSP_bh34_ch2_0(30); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w4_1 <= DSP_bh34_ch2_0(29); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w3_1 <= DSP_bh34_ch2_0(28); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w2_1 <= DSP_bh34_ch2_0(27); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w1_1 <= DSP_bh34_ch2_0(26); -- cycle= 0 cp= 1.638e-09
   heap_bh34_w0_1 <= DSP_bh34_ch2_0(25); -- cycle= 0 cp= 1.638e-09
   ----------------Synchro barrier, entering cycle 0----------------

   -- Adding the constant bits
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   finalAdderIn0_bh34 <= "0" & heap_bh34_w63_0_d1 & heap_bh34_w62_0_d1 & heap_bh34_w61_0_d1 & heap_bh34_w60_0_d1 & heap_bh34_w59_0_d1 & heap_bh34_w58_0_d1 & heap_bh34_w57_0_d1 & heap_bh34_w56_0_d1 & heap_bh34_w55_0_d1 & heap_bh34_w54_0_d1 & heap_bh34_w53_0_d1 & heap_bh34_w52_0_d1 & heap_bh34_w51_0_d1 & heap_bh34_w50_0_d1 & heap_bh34_w49_0_d1 & heap_bh34_w48_0_d1 & heap_bh34_w47_0_d1 & heap_bh34_w46_0_d1 & heap_bh34_w45_0_d1 & heap_bh34_w44_0_d1 & heap_bh34_w43_0_d1 & heap_bh34_w42_0_d1 & heap_bh34_w41_0_d1 & heap_bh34_w40_0_d1 & heap_bh34_w39_1_d1 & heap_bh34_w38_1_d1 & heap_bh34_w37_1_d1 & heap_bh34_w36_1_d1 & heap_bh34_w35_1_d1 & heap_bh34_w34_1_d1 & heap_bh34_w33_1_d1 & heap_bh34_w32_1_d1 & heap_bh34_w31_1_d1 & heap_bh34_w30_1_d1 & heap_bh34_w29_1_d1 & heap_bh34_w28_1_d1 & heap_bh34_w27_1_d1 & heap_bh34_w26_1_d1 & heap_bh34_w25_1_d1 & heap_bh34_w24_1_d1 & heap_bh34_w23_1_d1 & heap_bh34_w22_0_d1 & heap_bh34_w21_0_d1 & heap_bh34_w20_0_d1 & heap_bh34_w19_0_d1 & heap_bh34_w18_0_d1 & heap_bh34_w17_0_d1 & heap_bh34_w16_0_d1 & heap_bh34_w15_1_d1 & heap_bh34_w14_1_d1 & heap_bh34_w13_1_d1 & heap_bh34_w12_1_d1 & heap_bh34_w11_1_d1 & heap_bh34_w10_1_d1 & heap_bh34_w9_1_d1 & heap_bh34_w8_1_d1 & heap_bh34_w7_1_d1 & heap_bh34_w6_1_d1 & heap_bh34_w5_1_d1 & heap_bh34_w4_1_d1 & heap_bh34_w3_1_d1 & heap_bh34_w2_1_d1 & heap_bh34_w1_1_d1 & heap_bh34_w0_1_d1;
   finalAdderIn1_bh34 <= "0" & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh34_w39_0_d1 & heap_bh34_w38_0_d1 & heap_bh34_w37_0_d1 & heap_bh34_w36_0_d1 & heap_bh34_w35_0_d1 & heap_bh34_w34_0_d1 & heap_bh34_w33_0_d1 & heap_bh34_w32_0_d1 & heap_bh34_w31_0_d1 & heap_bh34_w30_0_d1 & heap_bh34_w29_0_d1 & heap_bh34_w28_0_d1 & heap_bh34_w27_0_d1 & heap_bh34_w26_0_d1 & heap_bh34_w25_0_d1 & heap_bh34_w24_0_d1 & heap_bh34_w23_0_d1 & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh34_w15_0_d1 & heap_bh34_w14_0_d1 & heap_bh34_w13_0_d1 & heap_bh34_w12_0_d1 & heap_bh34_w11_0_d1 & heap_bh34_w10_0_d1 & heap_bh34_w9_0_d1 & heap_bh34_w8_0_d1 & heap_bh34_w7_0_d1 & heap_bh34_w6_0_d1 & heap_bh34_w5_0_d1 & heap_bh34_w4_0_d1 & heap_bh34_w3_0_d1 & heap_bh34_w2_0_d1 & heap_bh34_w1_0_d1 & heap_bh34_w0_0_d1;
   finalAdderCin_bh34 <= '0';
   Adder_final34_0: IntAdder_65_f400_uid45  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => finalAdderCin_bh34,
                 R => finalAdderOut_bh34   ,
                 X => finalAdderIn0_bh34,
                 Y => finalAdderIn1_bh34);
   -- concatenate all the compressed chunks
   CompressionResult34 <= finalAdderOut_bh34;
   -- End of code generated by BitHeap::generateCompressorVHDL
   R <= CompressionResult34(63 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_66_f400_uid53
--                     (IntAdderClassical_66_f400_uid55)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_66_f400_uid53 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(65 downto 0);
          Y : in  std_logic_vector(65 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(65 downto 0)   );
end entity;

architecture arch of IntAdder_66_f400_uid53 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_66_f400_uid60
--                     (IntAdderClassical_66_f400_uid62)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_66_f400_uid60 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(65 downto 0);
          Y : in  std_logic_vector(65 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(65 downto 0)   );
end entity;

architecture arch of IntAdder_66_f400_uid60 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_61_f400_uid80
--                     (IntAdderClassical_61_f400_uid82)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_61_f400_uid80 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(60 downto 0);
          Y : in  std_logic_vector(60 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(60 downto 0)   );
end entity;

architecture arch of IntAdder_61_f400_uid80 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               IntMultiplier_UsingDSP_11_49_0_unsigned_uid67
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_11_49_0_unsigned_uid67 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          Y : in  std_logic_vector(48 downto 0);
          R : out  std_logic_vector(59 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_11_49_0_unsigned_uid67 is
   component IntAdder_61_f400_uid80 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(60 downto 0);
             Y : in  std_logic_vector(60 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(60 downto 0)   );
   end component;

signal XX_m68 :  std_logic_vector(48 downto 0);
signal YY_m68 :  std_logic_vector(10 downto 0);
signal DSP_bh69_ch0_0 :  std_logic_vector(40 downto 0);
signal heap_bh69_w59_0, heap_bh69_w59_0_d1 : std_logic;
signal heap_bh69_w58_0, heap_bh69_w58_0_d1 : std_logic;
signal heap_bh69_w57_0, heap_bh69_w57_0_d1 : std_logic;
signal heap_bh69_w56_0, heap_bh69_w56_0_d1 : std_logic;
signal heap_bh69_w55_0, heap_bh69_w55_0_d1 : std_logic;
signal heap_bh69_w54_0, heap_bh69_w54_0_d1 : std_logic;
signal heap_bh69_w53_0, heap_bh69_w53_0_d1 : std_logic;
signal heap_bh69_w52_0, heap_bh69_w52_0_d1 : std_logic;
signal heap_bh69_w51_0, heap_bh69_w51_0_d1 : std_logic;
signal heap_bh69_w50_0, heap_bh69_w50_0_d1 : std_logic;
signal heap_bh69_w49_0, heap_bh69_w49_0_d1 : std_logic;
signal heap_bh69_w48_0, heap_bh69_w48_0_d1 : std_logic;
signal heap_bh69_w47_0, heap_bh69_w47_0_d1 : std_logic;
signal heap_bh69_w46_0, heap_bh69_w46_0_d1 : std_logic;
signal heap_bh69_w45_0, heap_bh69_w45_0_d1 : std_logic;
signal heap_bh69_w44_0, heap_bh69_w44_0_d1 : std_logic;
signal heap_bh69_w43_0, heap_bh69_w43_0_d1 : std_logic;
signal heap_bh69_w42_0, heap_bh69_w42_0_d1 : std_logic;
signal heap_bh69_w41_0, heap_bh69_w41_0_d1 : std_logic;
signal heap_bh69_w40_0, heap_bh69_w40_0_d1 : std_logic;
signal heap_bh69_w39_0, heap_bh69_w39_0_d1 : std_logic;
signal heap_bh69_w38_0, heap_bh69_w38_0_d1 : std_logic;
signal heap_bh69_w37_0, heap_bh69_w37_0_d1 : std_logic;
signal heap_bh69_w36_0, heap_bh69_w36_0_d1 : std_logic;
signal heap_bh69_w35_0, heap_bh69_w35_0_d1 : std_logic;
signal heap_bh69_w34_0, heap_bh69_w34_0_d1 : std_logic;
signal heap_bh69_w33_0, heap_bh69_w33_0_d1 : std_logic;
signal heap_bh69_w32_0, heap_bh69_w32_0_d1 : std_logic;
signal heap_bh69_w31_0, heap_bh69_w31_0_d1 : std_logic;
signal heap_bh69_w30_0, heap_bh69_w30_0_d1 : std_logic;
signal heap_bh69_w29_0, heap_bh69_w29_0_d1 : std_logic;
signal heap_bh69_w28_0, heap_bh69_w28_0_d1 : std_logic;
signal heap_bh69_w27_0, heap_bh69_w27_0_d1 : std_logic;
signal heap_bh69_w26_0, heap_bh69_w26_0_d1 : std_logic;
signal heap_bh69_w25_0, heap_bh69_w25_0_d1 : std_logic;
signal heap_bh69_w24_0, heap_bh69_w24_0_d1 : std_logic;
signal heap_bh69_w23_0, heap_bh69_w23_0_d1 : std_logic;
signal heap_bh69_w22_0, heap_bh69_w22_0_d1 : std_logic;
signal heap_bh69_w21_0, heap_bh69_w21_0_d1 : std_logic;
signal heap_bh69_w20_0, heap_bh69_w20_0_d1 : std_logic;
signal heap_bh69_w19_0, heap_bh69_w19_0_d1 : std_logic;
signal DSP_bh69_ch1_0 :  std_logic_vector(40 downto 0);
signal heap_bh69_w35_1, heap_bh69_w35_1_d1 : std_logic;
signal heap_bh69_w34_1, heap_bh69_w34_1_d1 : std_logic;
signal heap_bh69_w33_1, heap_bh69_w33_1_d1 : std_logic;
signal heap_bh69_w32_1, heap_bh69_w32_1_d1 : std_logic;
signal heap_bh69_w31_1, heap_bh69_w31_1_d1 : std_logic;
signal heap_bh69_w30_1, heap_bh69_w30_1_d1 : std_logic;
signal heap_bh69_w29_1, heap_bh69_w29_1_d1 : std_logic;
signal heap_bh69_w28_1, heap_bh69_w28_1_d1 : std_logic;
signal heap_bh69_w27_1, heap_bh69_w27_1_d1 : std_logic;
signal heap_bh69_w26_1, heap_bh69_w26_1_d1 : std_logic;
signal heap_bh69_w25_1, heap_bh69_w25_1_d1 : std_logic;
signal heap_bh69_w24_1, heap_bh69_w24_1_d1 : std_logic;
signal heap_bh69_w23_1, heap_bh69_w23_1_d1 : std_logic;
signal heap_bh69_w22_1, heap_bh69_w22_1_d1 : std_logic;
signal heap_bh69_w21_1, heap_bh69_w21_1_d1 : std_logic;
signal heap_bh69_w20_1, heap_bh69_w20_1_d1 : std_logic;
signal heap_bh69_w19_1, heap_bh69_w19_1_d1 : std_logic;
signal heap_bh69_w18_0, heap_bh69_w18_0_d1 : std_logic;
signal heap_bh69_w17_0, heap_bh69_w17_0_d1 : std_logic;
signal heap_bh69_w16_0, heap_bh69_w16_0_d1 : std_logic;
signal heap_bh69_w15_0, heap_bh69_w15_0_d1 : std_logic;
signal heap_bh69_w14_0, heap_bh69_w14_0_d1 : std_logic;
signal heap_bh69_w13_0, heap_bh69_w13_0_d1 : std_logic;
signal heap_bh69_w12_0, heap_bh69_w12_0_d1 : std_logic;
signal heap_bh69_w11_0, heap_bh69_w11_0_d1 : std_logic;
signal heap_bh69_w10_0, heap_bh69_w10_0_d1 : std_logic;
signal heap_bh69_w9_0, heap_bh69_w9_0_d1 : std_logic;
signal heap_bh69_w8_0, heap_bh69_w8_0_d1 : std_logic;
signal heap_bh69_w7_0, heap_bh69_w7_0_d1 : std_logic;
signal heap_bh69_w6_0, heap_bh69_w6_0_d1 : std_logic;
signal heap_bh69_w5_0, heap_bh69_w5_0_d1 : std_logic;
signal heap_bh69_w4_0, heap_bh69_w4_0_d1 : std_logic;
signal heap_bh69_w3_0, heap_bh69_w3_0_d1 : std_logic;
signal heap_bh69_w2_0, heap_bh69_w2_0_d1 : std_logic;
signal heap_bh69_w1_0, heap_bh69_w1_0_d1 : std_logic;
signal heap_bh69_w0_0, heap_bh69_w0_0_d1 : std_logic;
signal DSP_bh69_ch2_0 :  std_logic_vector(40 downto 0);
signal heap_bh69_w11_1, heap_bh69_w11_1_d1 : std_logic;
signal heap_bh69_w10_1, heap_bh69_w10_1_d1 : std_logic;
signal heap_bh69_w9_1, heap_bh69_w9_1_d1 : std_logic;
signal heap_bh69_w8_1, heap_bh69_w8_1_d1 : std_logic;
signal heap_bh69_w7_1, heap_bh69_w7_1_d1 : std_logic;
signal heap_bh69_w6_1, heap_bh69_w6_1_d1 : std_logic;
signal heap_bh69_w5_1, heap_bh69_w5_1_d1 : std_logic;
signal heap_bh69_w4_1, heap_bh69_w4_1_d1 : std_logic;
signal heap_bh69_w3_1, heap_bh69_w3_1_d1 : std_logic;
signal heap_bh69_w2_1, heap_bh69_w2_1_d1 : std_logic;
signal heap_bh69_w1_1, heap_bh69_w1_1_d1 : std_logic;
signal heap_bh69_w0_1, heap_bh69_w0_1_d1 : std_logic;
signal finalAdderIn0_bh69 :  std_logic_vector(60 downto 0);
signal finalAdderIn1_bh69 :  std_logic_vector(60 downto 0);
signal finalAdderCin_bh69 : std_logic;
signal finalAdderOut_bh69 :  std_logic_vector(60 downto 0);
signal CompressionResult69 :  std_logic_vector(60 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            heap_bh69_w59_0_d1 <=  heap_bh69_w59_0;
            heap_bh69_w58_0_d1 <=  heap_bh69_w58_0;
            heap_bh69_w57_0_d1 <=  heap_bh69_w57_0;
            heap_bh69_w56_0_d1 <=  heap_bh69_w56_0;
            heap_bh69_w55_0_d1 <=  heap_bh69_w55_0;
            heap_bh69_w54_0_d1 <=  heap_bh69_w54_0;
            heap_bh69_w53_0_d1 <=  heap_bh69_w53_0;
            heap_bh69_w52_0_d1 <=  heap_bh69_w52_0;
            heap_bh69_w51_0_d1 <=  heap_bh69_w51_0;
            heap_bh69_w50_0_d1 <=  heap_bh69_w50_0;
            heap_bh69_w49_0_d1 <=  heap_bh69_w49_0;
            heap_bh69_w48_0_d1 <=  heap_bh69_w48_0;
            heap_bh69_w47_0_d1 <=  heap_bh69_w47_0;
            heap_bh69_w46_0_d1 <=  heap_bh69_w46_0;
            heap_bh69_w45_0_d1 <=  heap_bh69_w45_0;
            heap_bh69_w44_0_d1 <=  heap_bh69_w44_0;
            heap_bh69_w43_0_d1 <=  heap_bh69_w43_0;
            heap_bh69_w42_0_d1 <=  heap_bh69_w42_0;
            heap_bh69_w41_0_d1 <=  heap_bh69_w41_0;
            heap_bh69_w40_0_d1 <=  heap_bh69_w40_0;
            heap_bh69_w39_0_d1 <=  heap_bh69_w39_0;
            heap_bh69_w38_0_d1 <=  heap_bh69_w38_0;
            heap_bh69_w37_0_d1 <=  heap_bh69_w37_0;
            heap_bh69_w36_0_d1 <=  heap_bh69_w36_0;
            heap_bh69_w35_0_d1 <=  heap_bh69_w35_0;
            heap_bh69_w34_0_d1 <=  heap_bh69_w34_0;
            heap_bh69_w33_0_d1 <=  heap_bh69_w33_0;
            heap_bh69_w32_0_d1 <=  heap_bh69_w32_0;
            heap_bh69_w31_0_d1 <=  heap_bh69_w31_0;
            heap_bh69_w30_0_d1 <=  heap_bh69_w30_0;
            heap_bh69_w29_0_d1 <=  heap_bh69_w29_0;
            heap_bh69_w28_0_d1 <=  heap_bh69_w28_0;
            heap_bh69_w27_0_d1 <=  heap_bh69_w27_0;
            heap_bh69_w26_0_d1 <=  heap_bh69_w26_0;
            heap_bh69_w25_0_d1 <=  heap_bh69_w25_0;
            heap_bh69_w24_0_d1 <=  heap_bh69_w24_0;
            heap_bh69_w23_0_d1 <=  heap_bh69_w23_0;
            heap_bh69_w22_0_d1 <=  heap_bh69_w22_0;
            heap_bh69_w21_0_d1 <=  heap_bh69_w21_0;
            heap_bh69_w20_0_d1 <=  heap_bh69_w20_0;
            heap_bh69_w19_0_d1 <=  heap_bh69_w19_0;
            heap_bh69_w35_1_d1 <=  heap_bh69_w35_1;
            heap_bh69_w34_1_d1 <=  heap_bh69_w34_1;
            heap_bh69_w33_1_d1 <=  heap_bh69_w33_1;
            heap_bh69_w32_1_d1 <=  heap_bh69_w32_1;
            heap_bh69_w31_1_d1 <=  heap_bh69_w31_1;
            heap_bh69_w30_1_d1 <=  heap_bh69_w30_1;
            heap_bh69_w29_1_d1 <=  heap_bh69_w29_1;
            heap_bh69_w28_1_d1 <=  heap_bh69_w28_1;
            heap_bh69_w27_1_d1 <=  heap_bh69_w27_1;
            heap_bh69_w26_1_d1 <=  heap_bh69_w26_1;
            heap_bh69_w25_1_d1 <=  heap_bh69_w25_1;
            heap_bh69_w24_1_d1 <=  heap_bh69_w24_1;
            heap_bh69_w23_1_d1 <=  heap_bh69_w23_1;
            heap_bh69_w22_1_d1 <=  heap_bh69_w22_1;
            heap_bh69_w21_1_d1 <=  heap_bh69_w21_1;
            heap_bh69_w20_1_d1 <=  heap_bh69_w20_1;
            heap_bh69_w19_1_d1 <=  heap_bh69_w19_1;
            heap_bh69_w18_0_d1 <=  heap_bh69_w18_0;
            heap_bh69_w17_0_d1 <=  heap_bh69_w17_0;
            heap_bh69_w16_0_d1 <=  heap_bh69_w16_0;
            heap_bh69_w15_0_d1 <=  heap_bh69_w15_0;
            heap_bh69_w14_0_d1 <=  heap_bh69_w14_0;
            heap_bh69_w13_0_d1 <=  heap_bh69_w13_0;
            heap_bh69_w12_0_d1 <=  heap_bh69_w12_0;
            heap_bh69_w11_0_d1 <=  heap_bh69_w11_0;
            heap_bh69_w10_0_d1 <=  heap_bh69_w10_0;
            heap_bh69_w9_0_d1 <=  heap_bh69_w9_0;
            heap_bh69_w8_0_d1 <=  heap_bh69_w8_0;
            heap_bh69_w7_0_d1 <=  heap_bh69_w7_0;
            heap_bh69_w6_0_d1 <=  heap_bh69_w6_0;
            heap_bh69_w5_0_d1 <=  heap_bh69_w5_0;
            heap_bh69_w4_0_d1 <=  heap_bh69_w4_0;
            heap_bh69_w3_0_d1 <=  heap_bh69_w3_0;
            heap_bh69_w2_0_d1 <=  heap_bh69_w2_0;
            heap_bh69_w1_0_d1 <=  heap_bh69_w1_0;
            heap_bh69_w0_0_d1 <=  heap_bh69_w0_0;
            heap_bh69_w11_1_d1 <=  heap_bh69_w11_1;
            heap_bh69_w10_1_d1 <=  heap_bh69_w10_1;
            heap_bh69_w9_1_d1 <=  heap_bh69_w9_1;
            heap_bh69_w8_1_d1 <=  heap_bh69_w8_1;
            heap_bh69_w7_1_d1 <=  heap_bh69_w7_1;
            heap_bh69_w6_1_d1 <=  heap_bh69_w6_1;
            heap_bh69_w5_1_d1 <=  heap_bh69_w5_1;
            heap_bh69_w4_1_d1 <=  heap_bh69_w4_1;
            heap_bh69_w3_1_d1 <=  heap_bh69_w3_1;
            heap_bh69_w2_1_d1 <=  heap_bh69_w2_1;
            heap_bh69_w1_1_d1 <=  heap_bh69_w1_1;
            heap_bh69_w0_1_d1 <=  heap_bh69_w0_1;
         end if;
      end process;
   XX_m68 <= Y ;
   YY_m68 <= X ;
   
   -- Beginning of code generated by BitHeap::generateCompressorVHDL
   -- code generated by BitHeap::generateSupertileVHDL()
   ----------------Synchro barrier, entering cycle 0----------------
   DSP_bh69_ch0_0 <= ("" & XX_m68(48 downto 25) & "") * ("" & YY_m68(10 downto 0) & "000000");
   heap_bh69_w59_0 <= DSP_bh69_ch0_0(40); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w58_0 <= DSP_bh69_ch0_0(39); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w57_0 <= DSP_bh69_ch0_0(38); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w56_0 <= DSP_bh69_ch0_0(37); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w55_0 <= DSP_bh69_ch0_0(36); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w54_0 <= DSP_bh69_ch0_0(35); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w53_0 <= DSP_bh69_ch0_0(34); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w52_0 <= DSP_bh69_ch0_0(33); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w51_0 <= DSP_bh69_ch0_0(32); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w50_0 <= DSP_bh69_ch0_0(31); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w49_0 <= DSP_bh69_ch0_0(30); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w48_0 <= DSP_bh69_ch0_0(29); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w47_0 <= DSP_bh69_ch0_0(28); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w46_0 <= DSP_bh69_ch0_0(27); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w45_0 <= DSP_bh69_ch0_0(26); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w44_0 <= DSP_bh69_ch0_0(25); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w43_0 <= DSP_bh69_ch0_0(24); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w42_0 <= DSP_bh69_ch0_0(23); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w41_0 <= DSP_bh69_ch0_0(22); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w40_0 <= DSP_bh69_ch0_0(21); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w39_0 <= DSP_bh69_ch0_0(20); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w38_0 <= DSP_bh69_ch0_0(19); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w37_0 <= DSP_bh69_ch0_0(18); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w36_0 <= DSP_bh69_ch0_0(17); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w35_0 <= DSP_bh69_ch0_0(16); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w34_0 <= DSP_bh69_ch0_0(15); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w33_0 <= DSP_bh69_ch0_0(14); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w32_0 <= DSP_bh69_ch0_0(13); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w31_0 <= DSP_bh69_ch0_0(12); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w30_0 <= DSP_bh69_ch0_0(11); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w29_0 <= DSP_bh69_ch0_0(10); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w28_0 <= DSP_bh69_ch0_0(9); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w27_0 <= DSP_bh69_ch0_0(8); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w26_0 <= DSP_bh69_ch0_0(7); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w25_0 <= DSP_bh69_ch0_0(6); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w24_0 <= DSP_bh69_ch0_0(5); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w23_0 <= DSP_bh69_ch0_0(4); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w22_0 <= DSP_bh69_ch0_0(3); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w21_0 <= DSP_bh69_ch0_0(2); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w20_0 <= DSP_bh69_ch0_0(1); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w19_0 <= DSP_bh69_ch0_0(0); -- cycle= 0 cp= 1.638e-09
   ----------------Synchro barrier, entering cycle 0----------------
   DSP_bh69_ch1_0 <= ("" & XX_m68(24 downto 1) & "") * ("" & YY_m68(10 downto 0) & "000000");
   heap_bh69_w35_1 <= DSP_bh69_ch1_0(40); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w34_1 <= DSP_bh69_ch1_0(39); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w33_1 <= DSP_bh69_ch1_0(38); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w32_1 <= DSP_bh69_ch1_0(37); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w31_1 <= DSP_bh69_ch1_0(36); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w30_1 <= DSP_bh69_ch1_0(35); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w29_1 <= DSP_bh69_ch1_0(34); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w28_1 <= DSP_bh69_ch1_0(33); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w27_1 <= DSP_bh69_ch1_0(32); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w26_1 <= DSP_bh69_ch1_0(31); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w25_1 <= DSP_bh69_ch1_0(30); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w24_1 <= DSP_bh69_ch1_0(29); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w23_1 <= DSP_bh69_ch1_0(28); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w22_1 <= DSP_bh69_ch1_0(27); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w21_1 <= DSP_bh69_ch1_0(26); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w20_1 <= DSP_bh69_ch1_0(25); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w19_1 <= DSP_bh69_ch1_0(24); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w18_0 <= DSP_bh69_ch1_0(23); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w17_0 <= DSP_bh69_ch1_0(22); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w16_0 <= DSP_bh69_ch1_0(21); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w15_0 <= DSP_bh69_ch1_0(20); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w14_0 <= DSP_bh69_ch1_0(19); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w13_0 <= DSP_bh69_ch1_0(18); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w12_0 <= DSP_bh69_ch1_0(17); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w11_0 <= DSP_bh69_ch1_0(16); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w10_0 <= DSP_bh69_ch1_0(15); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w9_0 <= DSP_bh69_ch1_0(14); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w8_0 <= DSP_bh69_ch1_0(13); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w7_0 <= DSP_bh69_ch1_0(12); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w6_0 <= DSP_bh69_ch1_0(11); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w5_0 <= DSP_bh69_ch1_0(10); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w4_0 <= DSP_bh69_ch1_0(9); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w3_0 <= DSP_bh69_ch1_0(8); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w2_0 <= DSP_bh69_ch1_0(7); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w1_0 <= DSP_bh69_ch1_0(6); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w0_0 <= DSP_bh69_ch1_0(5); -- cycle= 0 cp= 1.638e-09
   ----------------Synchro barrier, entering cycle 0----------------
   DSP_bh69_ch2_0 <= ("" & XX_m68(0 downto 0) & "00000000000000000000000") * ("" & YY_m68(10 downto 0) & "000000");
   heap_bh69_w11_1 <= DSP_bh69_ch2_0(40); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w10_1 <= DSP_bh69_ch2_0(39); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w9_1 <= DSP_bh69_ch2_0(38); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w8_1 <= DSP_bh69_ch2_0(37); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w7_1 <= DSP_bh69_ch2_0(36); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w6_1 <= DSP_bh69_ch2_0(35); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w5_1 <= DSP_bh69_ch2_0(34); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w4_1 <= DSP_bh69_ch2_0(33); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w3_1 <= DSP_bh69_ch2_0(32); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w2_1 <= DSP_bh69_ch2_0(31); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w1_1 <= DSP_bh69_ch2_0(30); -- cycle= 0 cp= 1.638e-09
   heap_bh69_w0_1 <= DSP_bh69_ch2_0(29); -- cycle= 0 cp= 1.638e-09
   ----------------Synchro barrier, entering cycle 0----------------

   -- Adding the constant bits
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   finalAdderIn0_bh69 <= "0" & heap_bh69_w59_0_d1 & heap_bh69_w58_0_d1 & heap_bh69_w57_0_d1 & heap_bh69_w56_0_d1 & heap_bh69_w55_0_d1 & heap_bh69_w54_0_d1 & heap_bh69_w53_0_d1 & heap_bh69_w52_0_d1 & heap_bh69_w51_0_d1 & heap_bh69_w50_0_d1 & heap_bh69_w49_0_d1 & heap_bh69_w48_0_d1 & heap_bh69_w47_0_d1 & heap_bh69_w46_0_d1 & heap_bh69_w45_0_d1 & heap_bh69_w44_0_d1 & heap_bh69_w43_0_d1 & heap_bh69_w42_0_d1 & heap_bh69_w41_0_d1 & heap_bh69_w40_0_d1 & heap_bh69_w39_0_d1 & heap_bh69_w38_0_d1 & heap_bh69_w37_0_d1 & heap_bh69_w36_0_d1 & heap_bh69_w35_1_d1 & heap_bh69_w34_1_d1 & heap_bh69_w33_1_d1 & heap_bh69_w32_1_d1 & heap_bh69_w31_1_d1 & heap_bh69_w30_1_d1 & heap_bh69_w29_1_d1 & heap_bh69_w28_1_d1 & heap_bh69_w27_1_d1 & heap_bh69_w26_1_d1 & heap_bh69_w25_1_d1 & heap_bh69_w24_1_d1 & heap_bh69_w23_1_d1 & heap_bh69_w22_1_d1 & heap_bh69_w21_1_d1 & heap_bh69_w20_1_d1 & heap_bh69_w19_1_d1 & heap_bh69_w18_0_d1 & heap_bh69_w17_0_d1 & heap_bh69_w16_0_d1 & heap_bh69_w15_0_d1 & heap_bh69_w14_0_d1 & heap_bh69_w13_0_d1 & heap_bh69_w12_0_d1 & heap_bh69_w11_1_d1 & heap_bh69_w10_1_d1 & heap_bh69_w9_1_d1 & heap_bh69_w8_1_d1 & heap_bh69_w7_1_d1 & heap_bh69_w6_1_d1 & heap_bh69_w5_1_d1 & heap_bh69_w4_1_d1 & heap_bh69_w3_1_d1 & heap_bh69_w2_1_d1 & heap_bh69_w1_1_d1 & heap_bh69_w0_1_d1;
   finalAdderIn1_bh69 <= "0" & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh69_w35_0_d1 & heap_bh69_w34_0_d1 & heap_bh69_w33_0_d1 & heap_bh69_w32_0_d1 & heap_bh69_w31_0_d1 & heap_bh69_w30_0_d1 & heap_bh69_w29_0_d1 & heap_bh69_w28_0_d1 & heap_bh69_w27_0_d1 & heap_bh69_w26_0_d1 & heap_bh69_w25_0_d1 & heap_bh69_w24_0_d1 & heap_bh69_w23_0_d1 & heap_bh69_w22_0_d1 & heap_bh69_w21_0_d1 & heap_bh69_w20_0_d1 & heap_bh69_w19_0_d1 & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh69_w11_0_d1 & heap_bh69_w10_0_d1 & heap_bh69_w9_0_d1 & heap_bh69_w8_0_d1 & heap_bh69_w7_0_d1 & heap_bh69_w6_0_d1 & heap_bh69_w5_0_d1 & heap_bh69_w4_0_d1 & heap_bh69_w3_0_d1 & heap_bh69_w2_0_d1 & heap_bh69_w1_0_d1 & heap_bh69_w0_0_d1;
   finalAdderCin_bh69 <= '0';
   Adder_final69_0: IntAdder_61_f400_uid80  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => finalAdderCin_bh69,
                 R => finalAdderOut_bh69   ,
                 X => finalAdderIn0_bh69,
                 Y => finalAdderIn1_bh69);
   -- concatenate all the compressed chunks
   CompressionResult69 <= finalAdderOut_bh69;
   -- End of code generated by BitHeap::generateCompressorVHDL
   R <= CompressionResult69(59 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_56_f400_uid88
--                     (IntAdderClassical_56_f400_uid90)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_56_f400_uid88 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(55 downto 0);
          Y : in  std_logic_vector(55 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntAdder_56_f400_uid88 is
signal X_d1 :  std_logic_vector(55 downto 0);
signal Y_d1 :  std_logic_vector(55 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
    R <= X_d1 + Y_d1 + Cin_d1;
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_56_f400_uid95
--                    (IntAdderAlternative_56_f400_uid99)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_56_f400_uid95 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(55 downto 0);
          Y : in  std_logic_vector(55 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntAdder_56_f400_uid95 is
signal s_sum_l0_idx0 :  std_logic_vector(52 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(4 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(51 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(3 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(4 downto 0);
signal sum_l1_idx1 :  std_logic_vector(3 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(51 downto 0)) + ( "0" & Y(51 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(55 downto 52)) + ( "0" & Y(55 downto 52));
   sum_l0_idx0 <= s_sum_l0_idx0(51 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(52 downto 52);
   sum_l0_idx1 <= s_sum_l0_idx1(3 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(4 downto 4);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(3 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(4 downto 4);
   R <= sum_l1_idx1(3 downto 0) & sum_l0_idx0_d1(51 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                            IntSquarer_31_uid102
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2009)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee; 
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
library work;
entity IntSquarer_31_uid102 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(30 downto 0);
          R : out  std_logic_vector(61 downto 0)   );
end entity;

architecture arch of IntSquarer_31_uid102 is
signal x0_16, x0_16_d1 :  std_logic_vector(17 downto 0);
signal x17_32, x17_32_d1, x17_32_d2 :  std_logic_vector(17 downto 0);
signal x17_32_shr, x17_32_shr_d1 :  std_logic_vector(17 downto 0);
signal p0, p0_d1, p0_d2, p0_d3 :  std_logic_vector(35 downto 0);
signal p1_x2, p1_x2_d1 :  std_logic_vector(35 downto 0);
signal s1, s1_d1, s1_d2 :  std_logic_vector(35 downto 0);
signal p2, p2_d1 :  std_logic_vector(35 downto 0);
signal s2, s2_d1 :  std_logic_vector(35 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            x0_16_d1 <=  x0_16;
            x17_32_d1 <=  x17_32;
            x17_32_d2 <=  x17_32_d1;
            x17_32_shr_d1 <=  x17_32_shr;
            p0_d1 <=  p0;
            p0_d2 <=  p0_d1;
            p0_d3 <=  p0_d2;
            p1_x2_d1 <=  p1_x2;
            s1_d1 <=  s1;
            s1_d2 <=  s1_d1;
            p2_d1 <=  p2;
            s2_d1 <=  s2;
         end if;
      end process;
   x0_16 <= "0" & X(16 downto 0);
   x17_32 <= "00" & "00" & X(30 downto 17);
   x17_32_shr <= "0" & "00" & X(30 downto 17) & "0";
   ----------------Synchro barrier, entering cycle 1----------------
   p0 <= x0_16_d1 * x0_16_d1;
   p1_x2 <= x17_32_shr_d1 * x0_16_d1;
   ----------------Synchro barrier, entering cycle 2----------------
   s1 <= p1_x2_d1 + ( "00000000000000000" & p0_d1(35 downto 17));
   p2 <= x17_32_d2 * x17_32_d2;
   ----------------Synchro barrier, entering cycle 3----------------
   s2 <= p2_d1 + ( "00000000000000000" & s1_d1(35 downto 17));
   ----------------Synchro barrier, entering cycle 4----------------
   R <= s2_d1(27 downto 0) & s1_d2(16 downto 0) & p0_d3(16 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_56_f400_uid105
--                    (IntAdderAlternative_56_f400_uid109)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_56_f400_uid105 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(55 downto 0);
          Y : in  std_logic_vector(55 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntAdder_56_f400_uid105 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                              LogTable_0_11_83
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity LogTable_0_11_83 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          Y : out  std_logic_vector(82 downto 0)   );
end entity;

architecture arch of LogTable_0_11_83 is
   -- Build a 2-D array type for the RoM
   subtype word_t is std_logic_vector(82 downto 0);
   type memory_t is array(0 to 2047) of word_t;
   function init_rom
      return memory_t is 
      variable tmp : memory_t := (
   "11111111111111111011111111111111110000000000000000000000000000000000000000000000000",
   "11111111111111111011111111111111110000000000000000000000000000000000000000000000000",
   "00000000000111111100000111111111111010101010111010101011000100010001101110111100111",
   "00000000001111111100100000000001000101011001010101100010001001001100110101011111010",
   "00000000010111111101001000000100010000010100010001100001010100011001110011111001111",
   "00000000011111111110000000001010011011101010110001000100111011110011100000110011100",
   "00000000100111111111001000010100100111110001111000111001111000011011110110000100111",
   "00000000110000000000100000100011110101000100110000101110000000110100101101010011100",
   "00000000111000000010001000111001000100000100100100000000101010111110100110110001100",
   "00000001000000000100000001010101010101011000100010110011010101111110010110011000111",
   "00000001001000000110001001111001101001101110000010011010011011001011010010010001010",
   "00000001010000001000100010100111000001111000011110001110000111000111011111000001110",
   "00000001011000001011001011011110011110110001011000011011011010000011010110000100100",
   "00000001100000001110000100100001000001011000011010110101010000001110000010100101110",
   "00000001101000010001001101101111101010110011010111100101110001110100010010001101110",
   "00000001110000010100100111001011011100001110001001111111101010101110110110100111100",
   "00000001111000011000010000110101010110111010110111001111101010000010010101101101111",
   "00000010000000011100001010101110011100010001101111001110001001010001100110011000110",
   "00000010001000100000010100110111101101110001001101010000111011100100010111111101000",
   "00000010010000100100101111010010001100111101111000111101000100100011100011000100111",
   "00000010011000101001011001111110111011100010100110111000110111001100100010111010011",
   "00000010100000101110010100111110111011010000011001011101111100011101010101110100000",
   "00000010101000110011100000010011001101111110100001101011100001111010100101001001011",
   "00000010110000111000111011111100110101101010011111111000110000010001010100000111001",
   "00000010111000111110100111111100110100011000000100100111001001110101110101110011010",
   "00000011000001000100100100010100001100010001010001010101010001000001001011000101100",
   "00000011001001001010110001000011111111100110011001010001010110101110101001001101001",
   "00000011010001010001001110001101010000101110000010001100010000111011001010010010110",
   "00000011011001010111111011110001000010000101000101001100011001000111101001011101010",
   "00000011100001011110111001110000010110001110101111100000110011000000001100010000010",
   "00000011101001100110001000001100001111110100100011010100011011001001011011111000000",
   "00000011110001101101100111000101110001100110011000100001011101110101110000100101111",
   "00000011111001110101010110011101111110011010011101100100110110000011110010011010011",
   "00000100000001111101010110010101111001001101011000010001110100100111110010001110100",
   "00000100001010000101100110101110100101000010000110100101101111100001011111000010111",
   "00000100010010001110000111101001000101000001111111011011111001011111111011010100110",
   "00000100011010010110111001000110011100011100110011100001100001110100110110101010100",
   "00000100100010011111111011000111101110101000101110001001111100011001010000100100110",
   "00000100101010101001001101101101111111000010010110000010110010000100101001010011001",
   "00000100110010110010110000111010010001001100101110001000011001011000100110000100010",
   "00000100111010111100100100101101101000110001010110011010010111100010001110100000010",
   "00000101000011000110101001001001001001100000001100110000001001110011001001010000110",
   "00000101001011010000111110001101110111001111101101101101110111010011011110010100010",
   "00000101010011011011100011111100110101111100110101011001001011001110100101101100000",
   "00000101011011100110011010010111001001101011000000001110010111011100001001110000010",
   "00000101100011110001100001011101110110100100001011110101011111100111000100101011001",
   "00000101100011110001100001011101110110100100001011110101011111100111000100101011001",
   "00000101101011111100111001010010000000111000110111110111101100110100000000101111111",
   "00000101110100001000100001110100101101000000000110110100101001101001000011111110101",
   "00000101111100010100011011000110111111010111011110111000000110111000001111011011001",
   "00000110000100100000100101001001111100100011001010101111101000101110011011010011000",
   "00000110001100101100111111111110101001001101111010100000011100101000011001000111111",
   "00000110010100111001101011100110001010001001000100011101010111101111100101101101000",
   "00000110011101000110101000000001100100001100100101111100111110000000010100111000110",
   "00000110100101010011110101010001111100010111000100001111110001111011000001101001100",
   "00000110101101100001010011011000010111101101101101010110101101000010001101010000000",
   "00000110110101101111000010010101111011011100011000111001100001000110111000101100000",
   "00000110111101111101000010001011101100110101101000111101100010000101000011111110011",
   "00000111000110001011010010111010110001010010101010111100011000110001111111001111011",
   "00000111001110011001110100100100001110010011011000011010111110011101111001111010010",
   "00000111010110101000100111001001001001011110011000000000100001001010111100101110010",
   "00000111011110110111101010101010101000100000111110001101110000111010111011101000010",
   "00000111100111000110111111001001110001001111001110010100010101110101101101000100011",
   "00000111101111010110100100100111101001100011111011001110001111001001110100011110001",
   "00000111110111100110011011000101010111100000101000010101011011001001001110001110000",
   "00000111111111110110100010100100000001001101101010011011101000000011101011101100100",
   "00000111111111110110100010100100000001001101101010011011101000000011101011101100100",
   "00001000001000000110111011000100101100111010001000100010001110000000101110011110010",
   "00001000010000010111100100101000100000111011111100110010010001111010110010000000000",
   "00001000011000101000011111010000100011101111110101010100110001011101010011101001110",
   "00001000100000111001101010111101111011111001010101001010111000000111101001010010110",
   "00001000101001001011000111110001110000000010110101000110011101010110010110111110101",
   "00001000110001011100110101101101000110111101100100100010101011110100110100110011000",
   "00001000111001101110110100110001000111100001101010011100110001111000110110001110000",
   "00001001000010000001000100111110111000101110000110001100111011001010000100110001110",
   "00001001001010010011100110010111100001101000110000011111010011010111000000010000111",
   "00001001010010100110011000111100001001011110011100001101010010011001010111000011000",
   "00001001011010111001011100101101110111100010110111010110110001101011101001100010011",
   "00001001100011001100110001101101110011010000101011111011101010110001101100001100001",
   "00001001101011100000010111111101000100001001100000110101011111010101111011111001111",
   "00001001101011100000010111111101000100001001100000110101011111010101111011111001111",
   "00001001110011110100001111011100110001110101111010110001001010011101011001000010111",
   "00001001111100001000011000001110000100000101011101001000111011010011111101101110010",
   "00001010000100011100110010010010000010101110101010111110011001010011000100011011101",
   "00001010001100110001011101101001110101101111000111110100110001100100010100100001000",
   "00001010010101000110011010010110100101001011011000101011001110000010001010010101110",
   "00001010011101011011101000011001011001001111000100110111010101111000010001100010000",
   "00001010100101110001000111110011011010001100110110111111110111100101101000000000010",
   "00001010101110000110111000100101110000011110011101110111011100100010000000111011100",
   "00001010110110011100111010110001100100100100101101010111100110001000111111010001010",
   "00001010111110110011001110010111111111000111011111011011110100101011111111110110111",
   "00001011000111001001110011011010001000110101110100111100110111101101101011011111111",
   "00001011001111100000101001111001001010100101110110101100001000001000001001111100110",
   "00001011001111100000101001111001001010100101110110101100001000001000001001111100110",
   "00001011010111110111110001110110001101010100110110001111001100000000001111000101110",
   "00001011100000001111001011010010011010000111001110111011100100000111011100000001011",
   "00001011101000100110110110001110111010001000100110110010100011001110101110010001111",
   "00001011110000111110110010101100110110101011101111011101001111001011110111110001010",
   "00001011111001010111000000101101011001001010100111001000101011110011011010011101011",
   "00001100000001101111100000010001101011000110011001100010001111101001000011010111010",
   "00001100001010001000010001011010110110000111100000110100000010101000100000101100110",
   "00001100010010100001010100001010000011111101100110100001100110101000101111101001100",
   "00001100011010111010101000100000011110011111100100100100101001111011011110100000100",
   "00001100100011010100001110011111001111101011100110001010000011101011000000100010010",
   "00001100100011010100001110011111001111101011100110001010000011101011000000100010010",
   "00001100101011101110000110000111100001100111001000101110111010011000010001001011110",
   "00001100110100001000001111011010011110011110111100111101110100011011000100111011001",
   "00001100111100100010101010011001010000100111000111101100010010100110100110010001101",
   "00001101000100111101010111000101000010011011000010111000010100110011111110001000001",
   "00001101001101011000010101011110111110011101011110100110001000110101000110111000101",
   "00001101010101110011100101101000001111011000100001111110000011010001101010011101111",
   "00001101011110001111000111100001111111111101101100001010100010110000001011100101011",
   "00001101100110101010111011001101011011000101110101010110011101001101011011001111011",
   "00001101101111000111000000101011101011110001001111101011010111100011111011110110010",
   "00001101101111000111000000101011101011110001001111101011010111100011111011110110010",
   "00001101110111100011010111111101111101000111101000010000000111100101110011110011101",
   "00001110000000000000000001000101011010011000001000000111100000001010110001110111011",
   "00001110001000011100111100000011001110111001010101001111000111110100100110000101000",
   "00001110010000111010001000111000100110001001010011011110011001101011110010100111011",
   "00001110011001010111100111100110101011101101100101100101110000110110111000001010000",
   "00001110100001110101011000001110101011010011001110001101111110001110000010000111000",
   "00001110101010010011011010110001110000101110110000110111101000101101010111010110010",
   "00001110110010110001101111010001000111111100010010111010111000000111110100100111010",
   "00001110111011010000010101101101111100111111011100100111001010011100110110010011000",
   "00001110111011010000010101101101111100111111011100100111001010011100110110010011000",
   "00001111000011101111001110001001011100000011011010000011010011110010110111101100010",
   "00001111001100001110011000100100110001011010111100001101101000111000101110011000101",
   "00001111010100101101110101000001001001100000011001111100010100010000001000111000100",
   "00001111011101001101100011011111110000110101110000111101110110000011011000000110111",
   "00001111100101101101100100000001110100000100100110111001101110101000001011110100111",
   "00001111101110001101110110101000011111111110001010010001010011110010001010101010000",
   "00001111110110101110011011010101000001011011010011100000110000110110101110101100111",
   "00001111111111001111010010001000100101011100100110000000010001100100110000011100000",
   "00001111111111001111010010001000100101011100100110000000010001100100110000011100000",
   "00010000000111110000011011000100011001001010010001000101010111110010001001111011010",
   "00010000010000010001110110001001101001110100010001000100011100000001011100111100100",
   "00010000011000110011100011011001100100110010010000010010011001000001100111001010110",
   "00010000100001010101100010110101010111100011101000000110100010001010001111111101101",
   "00010000101001110111110100011110001111101111100001111100100100110110011011111100100",
   "00010000110010011010011000010101011011000100111000010110110101000000010010111010011",
   "00010000111010111101001110011100000111011010011000000000100100011111100101010011110",
   "00010000111010111101001110011100000111011010011000000000100100011111100101010011110",
   "00010001000011100000010110110011100010101110100000110000100101101101011110110101110",
   "00010001001100000011110001011100111011000111100110101011111001001111110100011110111",
   "00010001010100100111011110011001011110110011110011001000100110101101111100011111101",
   "00010001011101001011011101101010011100001001000101110001000000110001011111101110010",
   "00010001100101101111101111010001000001100101010101100110110100010101010011111001010",
   "00010001101110010100010011001110011101101110010010000110100011000100101111001100001",
   "00010001110110111001001001100011111111010001100100001011001001001101100101110111110",
   "00010001110110111001001001100011111111010001100100001011001001001101100101110111110",
   "00010001111111011110010010010010110101000100101111010001101110100111000011010011111",
   "00010010001000000011101101011100001110000101010010011101100011001111110000010000110",
   "00010010010000101001011011000001011001011000101001011100000111000101011000110010010",
   "00010010011001001111011011000011100110001100001101101001011101011000000100101111100",
   "00010010100001110101101101100100000011110101010111010100101011011011110110010110010",
   "00010010101010011100010010100100000001110001011110100100100010111010100010110001110",
   "00010010101010011100010010100100000001110001011110100100100010111010100010110001110",
   "00010010110011000011001010000100101111100101111100011100010111101000011001011001101",
   "00010010111011101010010100000111011101000000001100000001000000111101101110101111000",
   "00010011000100010001110000101101011001110101101011011110000110111000000000110010100",
   "00010011001100111001011111110111110110000011111101001011011010100100101010111111001",
   "00010011010101100001100001101000000001110000101000110010011010111000000000011010111",
   "00010011011110001001110101111111001101001001011100010100000100010010100011110010000",
   "00010011011110001001110101111111001101001001011100010100000100010010100011110010000",
   "00010011100110110010011100111110101000100100001101001110101100110111010100110011111",
   "00010011101111011011010110100111100100011110111001100100001011110101001011101101101",
   "00010011111000000100100010111011010001011111101001000000001101000101111011100001101",
   "00010100000000101110000001111011000000010100101101111110110000100101010101000000101",
   "00010100001001010111110011101000000001110100100110110010110101100010100100001100111",
   "00010100010010000001111000000011100110111101111110101101010001101110100011010010011",
   "00010100010010000001111000000011100110111101111110101101010001101110100011010010011",
   "00010100011010101100001111001111000000110111101111000011110100101001011110000111110",
   "00010100100011010110111001001011100000110001000000011000010110110010000010001100001",
   "00010100101100000001110101111010011000000001001011100000010100111000110111011111001",
   "00010100110100101101000101011100111000000111111010101100010111011010011111010000110",
   "00010100111101011000100111110100010010101101001010110000000110000010010110010000010",
   "00010101000110000100011101000001111001100001001100001010000111011001011000100101100",
   "00010101000110000100011101000001111001100001001100001010000111011001011000100101100",
   "00010101001110110000100101000110111110011100100100001100001101000010100110000011011",
   "00010101010111011101000000000100110011100000001110000011101011101000000110001010100",
   "00010101100000001001101101111100101010110101011100000001111111011011001011111001100",
   "00010101101000110110101110101111110110101101111000100101011101001001111001101011000",
   "00010101110001100100000010011111101001100011100111100010001111001100100110101010110",
   "00010101110001100100000010011111101001100011100111100010001111001100100110101010110",
   "00010101111010010001101001001101010101111001000111001011011111001110000111010001100",
   "00010110000010111111100010111010001110011001010001011100101100010000111010111011000",
   "00010110001011101101101111100111100101110111011101000011001101010100000010010100111",
   "00010110010100011100001111010110101111001111011110101000000000011010000001100110010",
   "00010110011101001011000010001000111101100101101001111001100110010100110010011101010",
   "00010110100101111010000111111111100100000110110010110110001010111000101011010000101",
   "00010110100101111010000111111111100100000110110010110110001010111000101011010000101",
   "00010110101110101001100000111011110110001000001110110101111001111001100000010001001",
   "00010110110111011001001100111111000111000111110101110101100000110100000101001000010",
   "00010111000000001001001100001010101010101100000011100000111101000110110101001101000",
   "00010111001000111001011110011111110100100011111000011110010111011100001001111111100",
   "00010111010001101010000011111111111000100110111011011001001011101001000111100001111",
   "00010111010001101010000011111111111000100110111011011001001011101001000111100001111",
   "00010111011010011010111100101100001010110101011010001101011101100011000111001110111",
   "00010111100011001100001000100101111111011000001011010011011010101111001010010110111",
   "00010111101011111101100111101110101010100000101110101011001001001101011101110100001",
   "00010111110100101111011010000111100000101001001111001000100011000011111001110000011",
   "00010111111101100001011111110001110110010100100011011111011111001010000111111101100",
   "00010111111101100001011111110001110110010100100011011111011111001010000111111101100",
   "00011000000110010011111000101111000000001110001111110000000110111001111100101110000",
   "00011000001111000110100101000000010011001010100110010011011001000110101110100010011",
   "00011000010111111001100100100111000100000110101001000111111001111110011001101001000",
   "00011000100000101100110111100100101000001000001010111110110000010110111100111001001",
   "00011000100000101100110111100100101000001000001010111110110000010110111100111001001",
   "00011000101001100000011101111010010100011101110000101000110000001010111110011011111",
   "00011000110010010100010111101001011110011110110010000011110010001000000110111101000",
   "00011000111011001000100100110011011011101011011011101000011000110010000011001100000",
   "00011001000011111101000101011001100001101100101111010111100010111100111011111100000",
   "00011001001100110001111001011101000110010100100110001000101011100001110101011110101",
   "00011001001100110001111001011101000110010100100110001000101011100001110101011110101",
   "00011001010101100111000000111111011111011101110000110111110110110000000111111111000",
   "00011001011110011100011100000010000011001011111001110100001100111110100011001110000",
   "00011001100111010010001010100110000111101011100101101110100010111110110000011010001",
   "00011001110000001000001100101101000011010010010101001000001111110110000101111100100",
   "00011001111000111110100010011000001100011110100101100010010000011110100001001010001",
   "00011001111000111110100010011000001100011110100101100010010000011110100001001010001",
   "00011010000001110101001011101000111001110111110010101100011000110010011011001010011",
   "00011010001010101100001000100000100010001110010111110100110010100110001110011010111",
   "00011010010011100011011001000000011100011011110000110111101010010010100011010111100",
   "00011010011100011010111101001001111111100010011011101111001001010001111011001000000",
   "00011010011100011010111101001001111111100010011011101111001001010001111011001000000",
   "00011010100101010010110100111110100010101101111001100011011110010100110000000010110",
   "00011010101110001011000000011111011101010010101111111011010011101110100100011110101",
   "00011010110111000011011111101110000110101110101010001100010011011111011000111100111",
   "00011010111111111100010010101011110110101000011010101011111001011100000011011111110",
   "00011010111111111100010010101011110110101000011010101011111001011100000011011111110",
   "00011011001000110101011001011010000100101111111100000000010011011000100010101111011",
   "00011011010001101110110011111010001000111110010010010001101111010111000111111101001",
   "00011011011010101000100010001101011011010101101100011011110111111111010100000010001",
   "00011011100011100010100100010101010100000001100101011111011110111111100100000100100",
   "00011011101100011100111010010011001011010110100101110100010101111100101010111010011",
   "00011011101100011100111010010011001011010110100101110100010101111100101010111010011",
   "00011011110101010111100100001000011001110010100100011011010101010001110101110100001",
   "00011011111110010010100001110110010111111100101000010000110001100100011011000001001",
   "00011100000111001101110011011110011110100101001001011110111111001110010001110100000",
   "00011100010000001001011001000010000110100101110010110001000100100001110100011001010",
   "00011100010000001001011001000010000110100101110010110001000100100001110100011001010",
   "00011100011001000101010010100010101001000001100010100101111010001010101100100000110",
   "00011100100010000001100000000001011111000100101100100011011010001110001100101101011",
   "00011100101010111110000001100000000010000100111010101001111101101110011000100111101",
   "00011100110011111010110110111111101011100001001110101000001000110010111111100111001",
   "00011100110011111010110110111111101011100001001110101000001000110010111111100111001",
   "00011100111100111000000000100001110101000010000011001110100101011011001101101110111",
   "00011101000101110101011110000111111000011001001101100100001100111011010111101111110",
   "00011101001110110011001111110011001111100001111110011010100000001001100111101101001",
   "00011101010111110001010101100101010100100001000011100010001110011100110000011000011",
   "00011101010111110001010101100101010100100001000011100010001110011100110000011000011",
   "00011101100000101111101111011111100001100100101001000000001011100000001110100000010",
   "00011101101001101110011101100011010001000100011010100010010100000000011111101001110",
   "00011101110010101101011111110001111101100001100100110101000001010010110111010010010",
   "00011101110010101101011111110001111101100001100100110101000001010010110111010010010",
   "00011101111011101100110110001101000001100110110110111000101011111011111011010001011",
   "00011110000100101100100000110101111000001000100011010111011101010111110010000000000",
   "00011110001101101100011111101101111100000100100001111011010000100111001100111011010",
   "00011110010110101100110010110110101000100010010000100100000010000100111011001101010",
   "00011110010110101100110010110110101000100010010000100100000010000100111011001101010",
   "00011110011111101101011010010001011000110010110100111110001110100110010000111000100",
   "00011110101000101110010101111111101000010000111101111001100001101010001111110010010",
   "00011110110001101111100110000010110010100001000100011111110010111010100000001100111",
   "00011110111010110001001010011100010011010001001101101100010011000001001000000111100",
   "00011110111010110001001010011100010011010001001101101100010011000001001000000111100",
   "00011111000011110011000011001101100110011001001011100011000111110110110000100111001",
   "00011111001100110101010000011000000111111010011110101000111000001100001001110100001",
   "00011111010101110111110001111101010100000000010111011010100110110010011110101010001",
   "00011111010101110111110001111101010100000000010111011010100110110010011110101010001",
   "00011111011110111010100111111110100110111111110111100101111101000101101010011010101",
   "00011111100111111101110010011101011101010111110011100001100101011100000010110110111",
   "00011111110001000001010001011011010011110000110011100101110100111110101010101100100",
   "00011111111010000101000100111001100110111101010101100101100101001101100000101111100",
   "00011111111010000101000100111001100110111101010101100101100101001101100000101111100",
   "00100000000011001001001100111001110011111001101110000111011101010011000001000110100",
   "00100000001100001101101001011101010111101100001001111111001011001010001110100000000",
   "00100000010101010010011010100101101111100100101111100111001100011010111010101011010",
   "00100000010101010010011010100101101111100100101111100111001100011010111010101011010",
   "00100000011110010111100000010100011000111101100000011010100111001111000101101010000",
   "00100000100111011100111010101010110001011010011010001111010011000101001100011110000",
   "00100000110000100010101001101010010110101001011000110000010001100010100000110100000",
   "00100000111001101000101101010100100110100010010110111000010111001001000011111100010",
   "00100000111001101000101101010100100110100010010110111000010111001001000011111100010",
   "00100001000010101111000101101010111111000111010000001101000100010100011111111011010",
   "00100001001011110101110010101110111110100100000010011001101110100001011011010011001",
   "00100001010100111100110100100010000011001110101110101010111001100010100011111100111",
   "00100001010100111100110100100010000011001110101110101010111001100010100011111100111",
   "00100001011110000100001011000101101011100111011011001010000001000111001110111101101",
   "00100001100111001011110110011011010110011000010100011001010010110110101011111111111",
   "00100001110000010011110110100100100010010101101110101111111000100011101011101011011",
   "00100001111001011100001011100010101110011110000111110110010010111011111001010001100",
   "00100001111001011100001011100010101110011110000111110110010010111011111001010001100",
   "00100010000010100100110101010111011001111010001000000011000100110110101000111010010",
   "00100010001011101101110100000100000011111100100011110111101111000110011100010110100",
   "00100010010100110111000111101010001100000010011101011101111100110001000001010110100",
   "00100010010100110111000111101010001100000010011101011101111100110001000001010110100",
   "00100010011110000000110000001011010001110011000110000101000000010001001101011000010",
   "00100010100111001010101101101000110100111111111111011111100001000110011011011111111",
   "00100010110000010101000000000100010101100100111101100001011010010101010010000000010",
   "00100010110000010101000000000100010101100100111101100001011010010101010010000000010",
   "00100010111001011111100111011111010011101000000111011110001001111100110110011000010",
   "00100011000010101010100011111011001111011001111001100111010001000100010110111101101",
   "00100011001011110101110101011001101001010101000110101011000101000100110010101111011",
   "00100011001011110101110101011001101001010101000110101011000101000100110010101111011",
   "00100011010101000001011011111100000001111110111001010011110001110010001000011100010",
   "00100011011110001101010111100011111010000110110101100110101100100111110111001010101",
   "00100011100111011001101000010010110010100110111010100011111000111100011011100110111",
   "00100011100111011001101000010010110010100110111010100011111000111100011011100110111",
   "00100011110000100110001110001010001100100011100011100101111101011111010101111000111",
   "00100011111001110011001001001011101001001011101010000010001011000101100100111110000",
   "00100100000011000000011001011000101001111000100110101000110100101000000101011101110",
   "00100100000011000000011001011000101001111000100110101000110100101000000101011101110",
   "00100100001100001101111110110010110000001110010011000101111000011000000010101111010",
   "00100100010101011011111001011011011101111011001011100001111010101100101001111100110",
   "00100100011110101010001001010100010100111000010000000011010010001110001111110101000",
   "00100100100111111000101110011110110111001001000110001111100101100010011010110001000",
   "00100100100111111000101110011110110111001001000110001111100101100010011010110001000",
   "00100100110001000111101000111100100110111011111010101101011010011101000011110110001",
   "00100100111010010110111000101111000110101001100010100110010110111010000010010110100",
   "00100101000011100110011101110111111000110101011101001001010011100011010110010011000",
   "00100101000011100110011101110111111000110101011101001001010011100011010110010011000",
   "00100101001100110110011000011000100000001101110101001101000000000111100111011100000",
   "00100101010110000110101000010010011111101011100010110010111001100100101111001110010",
   "00100101010110000110101000010010011111101011100010110010111001100100101111001110010",
   "00100101011111010111001101100111011010010010001100101010010010001010100101001000001",
   "00100101101000101000001000011000110011010000001001110011101011011001100101110000010",
   "00100101110001111001011000101000001101111110100011000100100010000001001110001000000",
   "00100101110001111001011000101000001101111110100011000100100010000001001110001000000",
   "00100101111011001010111110010111001110000001010100101011001100000010000101100001000",
   "00100110000100011100111001100111010111000111001111110011001000110111110001001101100",
   "00100110001101101111001010011010001101001001111100001001100011101110001110100101000",
   "00100110001101101111001010011010001101001001111100001001100011101110001110100101000",
   "00100110010111000001110000110001010100001101111001100010001000000110110000110010100",
   "00100110100000010100101100101110010000100010100001011100001000110000100000100110010",
   "00100110101001100111111110010010100110100010001000100111111000111000011101100100000",
   "00100110101001100111111110010010100110100010001000100111111000111000011101100100000",
   "00100110110010111011100101011111111010110010000000101100010111110101000001000110101",
   "00100110111100001111100010010111110010000010011001101101001111010001000100110100110",
   "00100111000101100011110100111011110001001110100011110001000011111010101110100011111",
   "00100111000101100011110100111011110001001110100011110001000011111010101110100011111",
   "00100111001110111000011101001101011101011100110000100111111000111001100101100111010",
   "00100111011000001101011011001110011011111110010101010010000101110000110101101100111",
   "00100111100001100010101111000000010010001111101011100111011111010001000101001010100",
   "00100111100001100010101111000000010010001111101011100111011111010001000101001010100",
   "00100111101010111000011000100100100101111000010011111110110010111110000101000010011",
   "00100111110100001110010111111100111100101010110110110101010101101100100010100110101",
   "00100111110100001110010111111100111100101010110110110101010101101100100010100110101",
   "00100111111101100100101101001010111100100101000110010111000100111100000011001010111",
   "00101000000110111011011000010000001011110000000000000110111011010001010011110001010",
   "00101000010000010010011001001110010000011111101110100111010111110100110111101001100",
   "00101000010000010010011001001110010000011111101110100111010111110100110111101001100",
   "00101000011001101001110000000110110001010011101011000011011000111010100001011001110",
   "00101000100011000001011100111011010100110110011110110111101001110101100011101110010",
   "00101000101100011001011111101101100001111110000101011100000011111110000111110010110",
   "00101000101100011001011111101101100001111110000101011100000011111110000111110010110",
   "00101000110101110001111000011110111111101011101101101101100011001011111000011011111",
   "00101000111111001010100111010001010101001011111011111000001101101010010010001111111",
   "00101001001000100011101100000110001001110110101011000001101111001010101001111110111",
   "00101001001000100011101100000110001001110110101011000001101111001010101001111110111",
   "00101001010001111101000110111111000101001111001110110100000111111000011011100101111",
   "00101001011011010110110111111101101111000100010101001000101110110011110101011011101",
   "00101001011011010110110111111101101111000100010101001000101110110011110101011011101",
   "00101001100100110000111111000011101111010000000111110011100111110111010100001101110",
   "00101001101110001011011100010010101101111000001110001111001101101100000101011100010",
   "00101001110111100110001111101100010011001101101111001000001111010010000111001000110",
   "00101001110111100110001111101100010011001101101111001000001111010010000111001000110",
   "00101010000001000001011001010010000111101101010010001010000001011111111100110110101",
   "00101010001010011100111001000101110011111111000001101011000100011110110011000000111",
   "00101010001010011100111001000101110011111111000001101011000100011110110011000000111",
   "00101010010011111000101111001001000000110110101100011001111101000111001010110100110",
   "00101010011101010100111011011101010111010011100111001010100010100010101010000111001",
   "00101010100110110001011110000100100000100000101110100011011111110111001011100100011",
   "00101010100110110001011110000100100000100000101110100011011111110111001011100100011",
   "00101010110000001110010111000000000101110100101000101100001010000000001101000100110",
   "00101010111001101011100110010001110000110001100110111010101001111010011010111000100",
   "00101010111001101011100110010001110000110001100110111010101001111010011010111000100",
   "00101011000011001001001011111011001011000101100111100010011011000110010111101000110",
   "00101011001100100111000111111101111110101010010111100010111110100110100010010110010",
   "00101011010110000101011010011011110101100101010100010111000010011101011100100111011",
   "00101011010110000101011010011011110101100101010100010111000010011101011100100111011",
   "00101011011111100100000011010110011010000111101101100011111101110000010100100101111",
   "00101011101001000011000010101111010110101110100110101001100001010010110111010011100",
   "00101011101001000011000010101111010110101110100110101001100001010010110111010011100",
   "00101011110010100010011000101000010110000010111000110001111101000000110001001101100",
   "00101011111100000010000101000011000010111001010100100010011010001001100011111111110",
   "00101100000101100010001000000001001000010010100011101011101010010011011001110111000",
   "00101100000101100010001000000001001000010010100011101011101010010011011001110111000",
   "00101100001111000010100001100100010001011011001010111011001011011001011111101100111",
   "00101100011000100011010001101110001001101011101011101100100000101010110000110111100",
   "00101100011000100011010001101110001001101011101011101100100000101010110000110111100",
   "00101100100010000100011000100000011100101000100101111011000000101101100000010100000",
   "00101100101011100101110101111100110110000010011001110011111000101100101100001111000",
   "00101100110101000111101010000101000001110101101001101000100100110011101010100000000",
   "00101100110101000111101010000101000001110101101001101000100100110011101010100000000",
   "00101100111110101001110100111010101100001010111011100001011101111100111101011001000",
   "00101101001000001100010110011111100001010110111011010000111100111001000001011011110",
   "00101101001000001100010110011111100001010110111011010000111100111001000001011011110",
   "00101101010001101111001110110101001101111010011100000110110010110001100110010101111",
   "00101101011011010010011101111101011110100010011010100011110111001110100110010011010",
   "00101101011011010010011101111101011110100010011010100011110111001110100110010011010",
   "00101101100100110110000011111010000000000111111110001110001100000001010000001001100",
   "00101101101110011010000000101100011111110000011011100101010110011010011010001101000",
   "00101101110111111110010100010110101010101101010101110111001110010000110100110010000",
   "00101101110111111110010100010110101010101101010101110111001110010000110100110010000",
   "00101110000001100010111110111010001110011100100000110101000010111100010100101111011",
   "00101110001011001000000000011000111000101000000010101000110110001010101111100111011",
   "00101110001011001000000000011000111000101000000010101000110110001010101111100111011",
   "00101110010100101101011000110100010111000110010101101011001100110011100100001111010",
   "00101110011110010011001000001110010111111010001010011001010101101111001100000000000",
   "00101110011110010011001000001110010111111010001010011001010101101111001100000000000",
   "00101110100111111001001110101000101001010010101001001011100110110110110010001110110",
   "00101110110001011111101100000100111001101011010100001100010000010001110000011101000",
   "00101110110001011111101100000100111001101011010100001100010000010001110000011101000",
   "00101110111011000110100000100100110111101100001001001110100101110101101111100100110",
   "00101111000100101101101100001010010010001001100011100110011110111110001111011011110",
   "00101111001110010101001110110110111000000100011110000000001101000000110111010111101",
   "00101111001110010101001110110110111000000100011110000000001101000000110111010111101",
   "00101111010111111101001000101100011000101010010100011000101000000011010011111001100",
   "00101111100001100101011001101100100011010101000101110101110010011000000110110100011",
   "00101111100001100101011001101100100011010101000101110101110010011000000110110100011",
   "00101111101011001110000001111001000111101011010110011111110010100111010000011110100",
   "00101111110100110111000001010011110101100000010001011010000100100111111010010000010",
   "00101111110100110111000001010011110101100000010001011010000100100111111010010000010",
   "00101111111110100000010111111110011100110011101010011101000001010000001011101010000",
   "00110000001000001010000101111010101101110010000000001111111101000000010100110011010",
   "00110000001000001010000101111010101101110010000000001111111101000000010100110011010",
   "00110000010001110100001011001010011000110100011110000011011101101110011010011000110",
   "00110000011011011110100111101111001110100000111101101100000111010111110000101101001",
   "00110000100101001001011011101010111111101010001001011101011111111101010100100000100",
   "00110000100101001001011011101010111111101010001001011101011111111101010100100000100",
   "00110000101110110100100110111111011101001111011110000101101010110000010010000011000",
   "00110000111000100000001001101110011000011101001100101000111010110100001011111001110",
   "00110000111000100000001001101110011000011101001100101000111010110100001011111001110",
   "00110001000010001100000011111001100010101100011100011101111100111011110100101010001",
   "00110001001011111000010101100010101101100011001101001010011001000110001111111001101",
   "00110001001011111000010101100010101101100011001101001010011001000110001111111001101",
   "00110001010101100100111110101011101010110100011000011111101011100001010000010111010",
   "00110001011111010001111111010110001100011111110100011000010101010110101010100010111",
   "00110001011111010001111111010110001100011111110100011000010101010110101010100010111",
   "00110001101000111111010111100100000100110010010100110101100101001001110100011101011",
   "00110001110010101101000111010111000110000101101101111101010111001010101100101101000",
   "00110001110010101101000111010111000110000101101101111101010111001010101100101101000",
   "00110001111100011011001110110001000011000000110101111000101101100100000100011000011",
   "00110010000110001001101101110011101110010111100110110010100000101010001000111001110",
   "00110010000110001001101101110011101110010111100110110010100000101010001000111001110",
   "00110010001111111000100100100000111011001011000000110110100111001111001100001010001",
   "00110010011001100111110010111010011100101001001100010001010111000011101010111101010",
   "00110010011001100111110010111010011100101001001100010001010111000011101010111101010",
   "00110010100011010111011001000010000110001101011011001111011101100111010011001010000",
   "00110010101101000111010110111001101011100000001011111110010001010000101100010100001",
   "00110010101101000111010110111001101011100000001011111110010001010000101100010100001",
   "00110010110110110111101100100011000000010111001010101100011010110001000111001111100",
   "00110011000000101000011001111111111000110101010011101010110111011001111010010000010",
   "00110011000000101000011001111111111000110101010011101010110111011001111010010000010",
   "00110011001010011001011111010010001001001010110101001110010011101001010001011110011",
   "00110011010100001010111100011011100101110101010001110000111110100011111011111110110",
   "00110011010100001010111100011011100101110101010001110000111110100011111011111110110",
   "00110011011101111100110001011110000011011111100001110100110110000001100000001001111",
   "00110011100111101110111110011011010111000001110110000110001011110001000011000100001",
   "00110011100111101110111110011011010111000001110110000110001011110001000011000100001",
   "00110011110001100001100011010101010101100001111001011110100011011011110000001111110",
   "00110011111011010100100000001101110100010010110011001000001001101011010000110010110",
   "00110011111011010100100000001101110100010010110011001000001001101011010000110010110",
   "00110100000101000111110101000110101000110101001000100001100100011001100010001011010",
   "00110100001110111011100010000001101000110110111111100001111100001111111110110000110",
   "00110100001110111011100010000001101000110110111111100001111100001111111110110000110",
   "00110100011000101111100111000000101010010100000000011101011111011011101011100110010",
   "00110100100010100100000100000101100011010101011000001010011101111100100000011111100",
   "00110100100010100100000100000101100011010101011000001010011101111100100000011111100",
   "00110100101100011000111001010010001010010001111010000110011111010101000001000101010",
   "00110100110110001110000110101000010101101110000010011100010010000000111111001000010",
   "00110100110110001110000110101000010101101110000010011100010010000000111111001000010",
   "00110101000000000011101100001001111100011011111000001001110100011000011111110010100",
   "00110101001001111001101001111000110101011011001111000110110111100101011111010101000",
   "00110101001001111001101001111000110101011011001111000110110111100101011111010101000",
   "00110101010011101111111111110110110111111001101010001011111100010001110000001101100",
   "00110101011101100110101110000101111011010010011101011001101001010011010100001110110",
   "00110101011101100110101110000101111011010010011101011001101001010011010100001110110",
   "00110101100111011101110100100111110111001110110000000000011100011101001111110011001",
   "00110101110001010101010011011110100011100101011110101000110101011010111001010101000",
   "00110101110001010101010011011110100011100101011110101000110101011010111001010101000",
   "00110101111011001101001010101011111000011011011101011011111010111011101000000100001",
   "00110110000101000101011010010001101110000011011010001100011010010101000111100011010",
   "00110110000101000101011010010001101110000011011010001100011010010101000111100011010",
   "00110110001110111110000010010001111100111101111110100000000001100010010110011000000",
   "00110110011000110111000010101110011101111001110001111001010011100101011000101010011",
   "00110110011000110111000010101110011101111001110001111001010011100101011000101010011",
   "00110110100010110000011011101001001001110011011100000001110111110010001000010011100",
   "00110110101100101010001101000011111001110101100110110101000011101000001110101010100",
   "00110110101100101010001101000011111001110101100110110101000011101000001110101010100",
   "00110110110110100100010111000000100111011001000000101010111111100010010101001000011",
   "00110111000000011110111001100001001100000100011110100100000110100000111011100111010",
   "00110111000000011110111001100001001100000100011110100100000110100000111011100111010",
   "00110111001010011001110100100111100001101100111110010101000000110111000101101101101",
   "00110111001010011001110100100111100001101100111110010101000000110111000101101101101",
   "00110111010100010101001000010101100010010101101000110010111001111111010001000100010",
   "00110111011110010000110100101101001000001111110100000000010001011110101000111111001",
   "00110111011110010000110100101101001000001111110100000000010001011110101000111111001",
   "00110111101000001100111001110000001101111011000101011010000111011101001101010110000",
   "00110111110010001001010111100000101110000101010100000101100100011001000100001111010",
   "00110111110010001001010111100000101110000101010100000101100100011001000100001111010",
   "00110111111100000110001110000000100011101010101010111101111100011011001111110111101",
   "00111000000110000011011101010001101001110101101011000011001110010100100011101000000",
   "00111000000110000011011101010001101001110101101011000011001110010100100011101000000",
   "00111000010000000001000101010101111011111111001101101000111110001000110101010001110",
   "00111000011001111111000110001111010101101110100110100101101011101111001000110111000",
   "00111000011001111111000110001111010101101110100110100101101011101111001000110111000",
   "00111000100011111101011111111111110010111001100110100010100101001101010111100100010",
   "00111000101101111100010010101001001111100100011101001011110101010101110011110110100",
   "00111000101101111100010010101001001111100100011101001011110101010101110011110110100",
   "00111000110111111011011110001101101000000001111011100001001110001101001110100110101",
   "00111000110111111011011110001101101000000001111011100001001110001101001110100110101",
   "00111001000001111011000010101110111000110011010110000111010000000000000011001001010",
   "00111001001011111011000000001110111110101000100111011000101100001101010001100011100",
   "00111001001011111011000000001110111110101000100111011000101100001101010001100011100",
   "00111001010101111011010110101111110110100000010001111000100101001101110000101000010",
   "00111001011111111100000110010011011101100111100010100100101010011110100010101010001",
   "00111001011111111100000110010011011101100111100010100100101010011110100010101010001",
   "00111001101001111101001110111011110001011010010011001000010001010100111001111100100",
   "00111001110011111110110000101010101111100011001100001111101010100010111011111011010",
   "00111001110011111110110000101010101111100011001100001111101010100010111011111011010",
   "00111001111110000000101011100010010101111011100111111011110100110011010011100000010",
   "00111001111110000000101011100010010101111011100111111011110100110011010011100000010",
   "00111010001000000010111111100100100010101011110011110110101100000011000101001001001",
   "00111010010010000101101100110011010100001010110011100111110110000000011001000100100",
   "00111010010010000101101100110011010100001010110011100111110110000000011001000100100",
   "00111010011100001000110011010000101000111110100011001001101011110100110001110110110",
   "00111010100110001100010010111110011111111011111000111111000001000010000111011111001",
   "00111010100110001100010010111110011111111011111000111111000001000010000111011111001",
   "00111010110000010000001011111110111000000110101000101001000111111001000000111110000",
   "00111010111010010100011110010011110000110001100100111110010011001111101000010111111",
   "00111010111010010100011110010011110000110001100100111110010011001111101000010111111",
   "00111011000100011001001001111111001001011110100010100000110101111111110111001011010",
   "00111011000100011001001001111111001001011110100010100000110101111111110111001011010",
   "00111011001110011110001111000011000001111110011001110110100000010011111010100111111",
   "00111011011000100011101101100001011010010001001010000000011010101000010001110101001",
   "00111011011000100011101101100001011010010001001010000000011010101000010001110101001",
   "00111011100010101001100101011100010010100101111010110011011110101010001001001110001",
   "00111011101100101111110110110101101011011010111111010001001110011001011000111000101",
   "00111011101100101111110110110101101011011010111111010001001110011001011000111000101",
   "00111011110110110110100001101111100101011101111000000001001001010101001101011001011",
   "00111011110110110110100001101111100101011101111000000001001001010101001101011001011",
   "00111100000000111101100110001100000001101011010101101010011111111010100100100011100",
   "00111100001011000101000100001101000001001111011011001110100101011011101001100100011",
   "00111100001011000101000100001101000001001111011011001110100101011011101001100100011",
   "00111100010101001100111011110100100101100101100000100011100000010111011110000111000",
   "00111100011111010101001101000100110000011000010100101111011001011000111111101110000",
   "00111100011111010101001101000100110000011000010100101111011001011000111111101110000",
   "00111100101001011101110111111111100011100010000000100100001001000100111011000000100",
   "00111100101001011101110111111111100011100010000000100100001001000100111011000000100",
   "00111100110011100110111100100111000001001100001000111011100100011101100000001010101",
   "00111100111101110000011010111101001011101111110001010100001000100011101110010000111",
   "00111100111101110000011010111101001011101111110001010100001000100011101110010000111",
   "00111101000111111010010011000100000101110101011110001110000100111101001100111001100",
   "00111101010010000100100100111101110010010101010111101001000101100110001101110011001",
   "00111101010010000100100100111101110010010101010111101001000101100110001101110011001",
   "00111101011100001111010000101100010100010111001011100010011011110111010010000000100",
   "00111101011100001111010000101100010100010111001011100010011011110111010010000000100",
   "00111101100110011010010110010001101111010010010000010011100111000101110000011000101",
   "00111101110000100101110101110000000110101101100111010001011100100110111101001101111",
   "00111101110000100101110101110000000110101101100111010001011100100110111101001101111",
   "00111101111010110001101111001001011110011111111111001011101111011101010100110100100",
   "00111101111010110001101111001001011110011111111111001011101111011101010100110100100",
   "00111110000100111110000010011111111010101111110110101101010111110111001101001000000",
   "00111110001111001010101111110101011111110011011110111100111010100110110100010011111",
   "00111110001111001010101111110101011111110011011110111100111010100110110100010011111",
   "00111110011001010111110111001100010010010000111101111101110000011011000100101111100",
   "00111110100011100101011000100110010110111110010001010001101101100000111000100000100",
   "00111110100011100101011000100110010110111110010001010001101101100000111000100000100",
   "00111110101101110011010100000101110011000001010000011011001001010100101001000011111",
   "00111110101101110011010100000101110011000001010000011011001001010100101001000011111",
   "00111110111000000001101001101100101011101111101111011111100110101011101001100110010",
   "00111111000010010000011001011101000110101111100001101010111100011101001100111101101",
   "00111111000010010000011001011101000110101111100001101010111100011101001100111101101",
   "00111111001100011111100011011001001001110110011011110010111110110011001010000011010",
   "00111111001100011111100011011001001001110110011011110010111110110011001010000011010",
   "00111111010110101111000111100010111011001010010110111011101001001001110011110110000",
   "00111111100000111111000101111100100001000001010010111011101001000110111100011101000",
   "00111111100000111111000101111100100001000001010010111011101001000110111100011101000",
   "00111111101011001111011110101000000010000001011001000001101010001111111100101100110",
   "00111111101011001111011110101000000010000001011001000001101010001111111100101100110",
   "00111111110101100000010001100111100101000000111110011010000011000110111100000000010",
   "00111111111111110001011110111101010001000110100110110101000011010110110110100101010",
   "00111111111111110001011110111101010001000110100110110101000011010110110110100101010",
   "01000000001010000011000110101011001101101001000111001101100011010110100010001011101",
   "01000000010100010101001000110011100010001111101000010000010101001010110011110110100",
   "01000000010100010101001000110011100010001111101000010000010101001010110011110110100",
   "01000000011110100111100101011000010110110001101001000011110111001111101011011110100",
   "01000000011110100111100101011000010110110001101001000011110111001111101011011110100",
   "01000000101000111010011100011011110011010111000001110000101000110000101100000110011",
   "01000000110011001101101110000000000000011000000110001001111111111000101010010110011",
   "01000000110011001101101110000000000000011000000110001001111111111000101010010110011",
   "01000000111101100001011010000111000110011101101000010111100010000000111100100011011",
   "01000000111101100001011010000111000110011101101000010111100010000000111100100011011",
   "01000001000111110101100000110011001110100000111011011110111110001000011010011100110",
   "01000001010010001010000010000110100001101011110110001110101001011010011100101111000",
   "01000001010010001010000010000110100001101011110110001110101001011010011100101111000",
   "01000001011100011110111110000011001001011000110101101000011110001110001110111110011",
   "01000001011100011110111110000011001001011000110101101000011110001110001110111110011",
   "01000001100110110100010100101011001111010010111111101101011101100110101000110100100",
   "01000001110001001010000110000000111101010110000110001001110011011011000101101110110",
   "01000001110001001010000110000000111101010110000110001001110011011011000101101110110",
   "01000001111011100000010010000110011101101110101001000001011101010001110100110111000",
   "01000001111011100000010010000110011101101110101001000001011101010001110100110111000",
   "01000010000101110110111000111101111010111001111001011101010100010011111101000110000",
   "01000010010000001101111010101001011111100101111100011000111010000011110011100111011",
   "01000010010000001101111010101001011111100101111100011000111010000011110011100111011",
   "01000010011010100101010111001011010110110001101101010000101000011110000101110011010",
   "01000010011010100101010111001011010110110001101101010000101000011110000101110011010",
   "01000010100100111101001110100101101011101101000000110000100101001110011001101001000",
   "01000010101111010101100000111010101001111000100111100011111000011111101010010100100",
   "01000010101111010101100000111010101001111000100111100011111000011111101010010100100",
   "01000010111001101110001110001100011101000110010001000100100111010001001001000001001",
   "01000010111001101110001110001100011101000110010001000100100111010001001001000001001",
   "01000011000100000111010110011101010001011000101110001100010001011000101100011110100",
   "01000011000100000111010110011101010001011000101110001100010001011000101100011110100",
   "01000011001110100000111001101111010011000011110100000100110011011010111100010001110",
   "01000011011000111010111000000100101110101100011110111010001100100010000111010101000",
   "01000011011000111010111000000100101110101100011110111010001100100010000111010101000",
   "01000011100011010101010001011111110001001000110100101100101000011100010111011110111",
   "01000011100011010101010001011111110001001000110100101100101000011100010111011110111",
   "01000011101101110000000110000010100111100000001000000011001101101010010110110000100",
   "01000011111000001011010101101111011111001010111010111111010000000110111101000111000",
   "01000011111000001011010101101111011111001010111010111111010000000110111101000111000",
   "01000100000010100111000000101000100101110011000001110000001000010001000000010000000",
   "01000100000010100111000000101000100101110011000001110000001000010001000000010000000",
   "01000100001101000011000110110000001001010011100101100111101111000000000001100100101",
   "01000100010111011111101000001000010111111001000111101111011110001100111000101101000",
   "01000100010111011111101000001000010111111001000111101111011110001100111000101101000",
   "01000100100001111100100100110011100000000001100011111101110110010111011011111010110",
   "01000100100001111100100100110011100000000001100011111101110110010111011011111010110",
   "01000100101100011001111100110011110000011100010011101100101001010010001010000100100",
   "01000100101100011001111100110011110000011100010011101100101001010010001010000100100",
   "01000100110110110111110000001011011000001010010000101111101001111100111100011010100",
   "01000101000001010101111110111100100110011101111000001100000001111000001001001101110",
   "01000101000001010101111110111100100110011101111000001100000001111000001001001101110",
   "01000101001011110100101001001001101010111011001101010000001011111001000010101101000",
   "01000101001011110100101001001001101010111011001101010000001011111001000010101101000",
   "01000101010110010011101110110100110101010111111100001100010100101001000000100100110",
   "01000101100000110011010000000000010101111011011101001011100000111000100100110010110",
   "01000101100000110011010000000000010101111011011101001011100000111000100100110010110",
   "01000101101011010011001100101110011100111110110111001101011001101111101111010010100",
   "01000101101011010011001100101110011100111110110111001101011001101111101111010010100",
   "01000101110101110011100101000001011011001101000011000000011111000100110110100101100",
   "01000101110101110011100101000001011011001101000011000000011111000100110110100101100",
   "01000110000000010100011000111011100001100010101101111101000000000011011110010010110",
   "01000110001010110101101000011111000001001110011101000000011010001100100110111110100",
   "01000110001010110101101000011111000001001110011101000000011010001100100110111110100",
   "01000110010101010111010011101110001011110000101111101001011110111001110101101000110",
   "01000110010101010111010011101110001011110000101111101001011110111001110101101000110",
   "01000110011111111001011010101011010010111100000010110100111111101100110011110110000",
   "01000110011111111001011010101011010010111100000010110100111111101100110011110110000",
   "01000110101010011011111101011000101000110100110011111011000001010100101100001011100",
   "01000110110100111110111011111000011111110001100011101100110101110011001001100011001",
   "01000110110100111110111011111000011111110001100011101100110101110011001001100011001",
   "01000110111111100010010110001101001010011010111001010011011101101010100010100011111",
   "01000110111111100010010110001101001010011010111001010011011101101010100010100011111",
   "01000111001010000110001100011000111011101011100101001110110000011110111101000010110",
   "01000111001010000110001100011000111011101011100101001110110000011110111101000010110",
   "01000111010100101010011110011110000110110000100100010101001100110011111000100001100",
   "01000111011111001111001100011110111111001001000010110100001111110000010001010110000",
   "01000111011111001111001100011110111111001001000010110100001111110000010001010110000",
   "01000111101001110100010110011101111000100110011111010001010100010010110000110111010",
   "01000111101001110100010110011101111000100110011111010001010100010010110000110111010",
   "01000111110100011001111100011101000111001100101101101011011010100000000010000110110",
   "01000111110100011001111100011101000111001100101101101011011010100000000010000110110",
   "01000111111110111111111110011110111111010001111010011101010110110101000101000000000",
   "01001000001001100110011100100101110101011110101101100000101001100111011101010011100",
   "01001000001001100110011100100101110101011110101101100000101001100111011101010011100",
   "01001000010100001101010110110011111110101110001101010000111110111101011101001000110",
   "01001000010100001101010110110011111110101110001101010000111110111101011101001000110",
   "01001000011110110100101101001011110000001110000001110000010111001000001101111100000",
   "01001000011110110100101101001011110000001110000001110000010111001000001101111100000",
   "01001000101001011100011111101111011111011110010111101011110111101001111101101010100",
   "01001000110100000100101110100001100010010010000011100001000101010010011000111001000",
   "01001000110100000100101110100001100010010010000011100001000101010010011000111001000",
   "01001000111110101101011001100100001110101110100100100100000110111011011101011101001",
   "01001000111110101101011001100100001110101110100100100100000110111011011101011101001",
   "01001001001001010110100000111001111011001100001000000110010001110000110100001111101",
   "01001001001001010110100000111001111011001100001000000110010001110000110100001111101",
   "01001001010100000000000100100100111110010101101100011101011110101100000011101111100",
   "01001001011110101010000100100111101111001001000100001100001001010000001111110111100",
   "01001001011110101010000100100111101111001001000100001100001001010000001111110111100",
   "01001001101001010100100001000100100100110110111001001001111000001110111110101101111",
   "01001001101001010100100001000100100100110110111001001001111000001110111110101101111",
   "01001001110011111111011001111101110111000010101111101100110000000001011100110101000",
   "01001001110011111111011001111101110111000010101111101100110000000001011100110101000",
   "01001001111110101010101111010101111101100011001001110011001110111111111110100101101",
   "01001001111110101010101111010101111101100011001001110011001110111111111110100101101",
   "01001010001001010110100001001111010000100001101010001110110100000010011111100001100",
   "01001010010100000010101111101100001000011010110111101111001111010100100011001111001",
   "01001010010100000010101111101100001000011010110111101111001111010100100011001111001",
   "01001010011110101111011010101110111101111110100000001110011101100111011110111000010",
   "01001010011110101111011010101110111101111110100000001110011101100111011110111000010",
   "01001010101001011100100010011010001010001111011011111101001110001101010101000110110",
   "01001010101001011100100010011010001010001111011011111101001110001101010101000110110",
   "01001010110100001010000110110000000110100011110000110000010011100111010001101000100",
   "01001010111110111000000111110011001100100100110101001110011111010010010100101000000",
   "01001010111110111000000111110011001100100100110101001110011111010010010100101000000",
   "01001011001001100110100101100101110110001111010011111111001000011101000001010011110",
   "01001011001001100110100101100101110110001111010011111111001000011101000001010011110",
   "01001011010100010101100000001010011101110011001110111001011110010001000110010101011",
   "01001011010100010101100000001010011101110011001110111001011110010001000110010101011",
   "01001011011111000100110111100011011101110100000010010100100101011011111001101100110",
   "01001011011111000100110111100011011101110100000010010100100101011011111001101100110",
   "01001011101001110100101011110011010001001000101000011000000001100000100101000110100",
   "01001011110100100100111100111100010010111011011100001101001001111111000010111110010",
   "01001011110100100100111100111100010010111011011100001101001001111111000010111110010",
   "01001011111111010101101011000000111110101010011101010001001011011010101111100001100",
   "01001011111111010101101011000000111110101010011101010001001011011010101111100001100",
   "01001100001010000110110110000011110000000111010010100111110100101100010100100001111",
   "01001100001010000110110110000011110000000111010010100111110100101100010100100001111",
   "01001100010100111000011110000111000011010111001110001110110000101001011001101111011",
   "01001100010100111000011110000111000011010111001110001110110000101001011001101111011",
   "01001100011111101010100011001101010100110011010000010001101100001101100111001011010",
   "01001100011111101010100011001101010100110011010000010001101100001101100111001011010",
   "01001100101010011101000101011001000001001000001010011111001001010000001001110011011",
   "01001100110101010000000100101100100101010110100011011101111110010001001110011110000",
   "01001100110101010000000100101100100101010110100011011101111110010001001110011110000",
   "01001101000000000011100001001010011110110010111010000011100011001010101010010001110",
   "01001101000000000011100001001010011110110010111010000011100011001010101010010001110",
   "01001101001010110111011010110101001011000101101000101010101011001111001010111110001",
   "01001101001010110111011010110101001011000101101000101010101011001111001010111110001",
   "01001101010101101011110001101111001000001011001000101011001100100011101101001101100",
   "01001101010101101011110001101111001000001011001000101011001100100011101101001101100",
   "01001101100000100000100101111010110100010011110101110010010100111110011010001001100",
   "01001101100000100000100101111010110100010011110101110010010100111110011010001001100",
   "01001101101011010101110111011010101110000100010001011011101100110110110000111100011",
   "01001101110110001011100110010001010100010101000110001011000111110010100100011101110",
   "01001101110110001011100110010001010100010101000110001011000111110010100100011101110",
   "01001110000001000001110010100001000110010011001011000111000011011011011000101111110",
   "01001110000001000001110010100001000110010011001011000111000011011011011000101111110",
   "01001110001011111000011100001100100011011111100111010011110100101000001111010010101",
   "01001110001011111000011100001100100011011111100111010011110100101000001111010010101",
   "01001110010110101111100011010110001011101111110101001111100011000111010100110011100",
   "01001110010110101111100011010110001011101111110101001111100011000111010100110011100",
   "01001110100001100111001000000000011111001101100110001110110011110011100110011010110",
   "01001110100001100111001000000000011111001101100110001110110011110011100110011010110",
   "01001110101100011111001010001101111110010111000101111010000010000010000111111110101",
   "01001110110111010111101010000001001001111110111101101011100111110011001000100101100",
   "01001110110111010111101010000001001001111110111101101011100111110011001000100101100",
   "01001111000010010000100111011100100011001100011000001110110101010010110110000001110",
   "01001111000010010000100111011100100011001100011000001110110101010010110110000001110",
   "01001111001101001010000010100010101011011011000100111111010111110110000011011001000",
   "01001111001101001010000010100010101011011011000100111111010111110110000011011001000",
   "01001111011000000011111011010110000100011011011011101001110000011110101010110001011",
   "01001111011000000011111011010110000100011011011011101001110000011110101010110001011",
   "01001111100010111110010001111001010000010010011111101100011010010100010101011111100",
   "01001111100010111110010001111001010000010010011111101100011010010100010101011111100",
   "01001111101101111001000110001110110001011010000011111001100000111101011010000000110",
   "01001111101101111001000110001110110001011010000011111001100000111101011010000000110",
   "01001111111000110100011000011001001010100000101101111001100111000100100010010011110",
   "01010000000011110000001000011010111110101001111001101110111101010111010001001000100",
   "01010000000011110000001000011010111110101001111001101110111101010111010001001000100",
   "01010000001110101100010110010110110001001101111101011001101010001010000000010111010",
   "01010000001110101100010110010110110001001101111101011001101010001010000000010111010",
   "01010000011001101001000010001111000101111010001100011100100001101101110110010010001",
   "01010000011001101001000010001111000101111010001100011100100001101101110110010010001",
   "01010000100100100110001100000110100000110000111011100010101111100100110011010111000",
   "01010000100100100110001100000110100000110000111011100010101111100100110011010111000",
   "01010000101111100011110011111111100110001001100100000110010001000000111101111101010",
   "01010000101111100011110011111111100110001001100100000110010001000000111101111101010",
   "01010000111010100001111001111100111010110000100111110111000000111011010101000001000",
   "01010000111010100001111001111100111010110000100111110111000000111011010101000001000",
   "01010001000101100000011110000001000011100111110100100010110101001110110110101101110",
   "01010001000101100000011110000001000011100111110100100010110101001110110110101101110",
   "01010001010000011111100000001110100110000110000111011110001110000100101011110010010",
   "01010001011011011111000000101000000111110111110001001101110110111110001100000110000",
   "01010001011011011111000000101000000111110111110001001101110110111110001100000110000",
   "01010001100110011110111111010000001110111110011001010000111010001001110100111010010",
   "01010001100110011110111111010000001110111110011001010000111010001001110100111010010",
   "01010001110001011111011100001001100001110001000001101100000110001111101101001100000",
   "01010001110001011111011100001001100001110001000001101100000110001111101101001100000",
   "01010001111100100000010111010110100110111100001010110101100110100010111000000001010",
   "01010001111100100000010111010110100110111100001010110101100110100010111000000001010",
   "01010010000111100001110000111010000101100001110111000001101110000100011001011101000",
   "01010010000111100001110000111010000101100001110111000001101110000100011001011101000",
   "01010010010010100011101000110110100100111001101110010000010101100101010101101100100",
   "01010010010010100011101000110110100100111001101110010000010101100101010101101100100",
   "01010010011101100101111111001110101100110001000001111011001100110100110110101111010",
   "01010010011101100101111111001110101100110001000001111011001100110100110110101111010",
   "01010010101000101000110100000101000101001010110000100100111111000111101000011011100",
   "01010010101000101000110100000101000101001010110000100100111111000111101000011011100",
   "01010010110011101100000111011100010110011111101001101001001011100101111110111110110",
   "01010010110011101100000111011100010110011111101001101001001011100101111110111110110",
   "01010010111110101111111001010111001001011110010001001100110001001101111111111101110",
   "01010011001001110100001001111000000111001011000011101111101110110111001001111010100",
   "01010011001001110100001001111000000111001011000011101111101110110111001001111010100",
   "01010011010100111000111001000001111001000000011001111111010111100100111010100111110",
   "01010011010100111000111001000001111001000000011001111111010111100100111010100111110",
   "01010011011111111110000110110111001000101110101100101001011011010101111000011011110",
   "01010011011111111110000110110111001000101110101100101001011011010101111000011011110",
   "01010011101011000011110011011010100000011100011000010000000100011101000110111001011",
   "01010011101011000011110011011010100000011100011000010000000100011101000110111001011",
   "01010011110110001001111110101110101010100110000000111110101001110011010011001110111",
   "01010011110110001001111110101110101010100110000000111110101001110011010011001110111",
   "01010100000001010000101000110110010001111110010110011111010110001101101001010100000",
   "01010100000001010000101000110110010001111110010110011111010110001101101001010100000",
   "01010100001100010111110001110100000001101110010111110001100101001000000101111101100",
   "01010100001100010111110001110100000001101110010111110001100101001000000101111101100",
   "01010100010111011111011001101010100101010101010111000001010100110000111111101001011",
   "01010100010111011111011001101010100101010101010111000001010100110000111111101001011",
   "01010100100010100111100000011100101000101000111101011111001110000100000010110010011",
   "01010100100010100111100000011100101000101000111101011111001110000100000010110010011",
   "01010100101101110000000110001100110111110101001111011001100010100010100011001110110",
   "01010100101101110000000110001100110111110101001111011001100010100010100011001110110",
   "01010100111000111001001010111101111111011100101111110110000000010111001000101010101",
   "01010100111000111001001010111101111111011100101111110110000000010111001000101010101",
   "01010101000100000010101110110010101100011000100100101100011100110011000000000100100",
   "01010101000100000010101110110010101100011000100100101100011100110011000000000100100",
   "01010101001111001100110001101101101011111000011010100010010101010011000000100100010",
   "01010101001111001100110001101101101011111000011010100010010101010011000000100100010",
   "01010101011010010111010011110001101011100010101000100111000111011010110110011111000",
   "01010101011010010111010011110001101011100010101000100111000111011010110110011111000",
   "01010101100101100010010101000001011001010100010100110001011111110100101011101011100",
   "01010101100101100010010101000001011001010100010100110001011111110100101011101011100",
   "01010101110000101101110101011111100011100001010111011101100000100011101000101001100",
   "01010101111011111001110101001110111000110100011111101011011110110111101110010111010",
   "01010101111011111001110101001110111000110100011111101011011110110111101110010111010",
   "01010110000111000110010100010010001000001111010110111111111000110001101101001001010",
   "01010110000111000110010100010010001000001111010110111111111000110001101101001001010",
   "01010110010010010011010010101100000001001010100101100100000010100101100001011010100",
   "01010110010010010011010010101100000001001010100101100100000010100101100001011010100",
   "01010110011101100000110000011111010011010101110110000111101100101010000011101001000",
   "01010110011101100000110000011111010011010101110110000111101100101010000011101001000",
   "01010110101000101110101101101110101110110111111010000011100001100100111101010000100",
   "01010110101000101110101101101110101110110111111010000011100001100100111101010000100",
   "01010110110011111101001010011101000100001110101101011100011101000001011000111100110",
   "01010110110011111101001010011101000100001110101101011100011101000001011000111100110",
   "01010110111111001100000110101101000100001111011011000111111011100000101001001011110",
   "01010110111111001100000110101101000100001111011011000111111011100000101001001011110",
   "01010111001010011011100010100001100000000110100000110001000011010011100100100000000",
   "01010111001010011011100010100001100000000110100000110001000011010011100100100000000",
   "01010111010101101011011101111101001001010111110010111110100110101011111011101011100",
   "01010111010101101011011101111101001001010111110010111110100110101011111011101011100",
   "01010111100000111011111001000010110001111110100001011001111111110100110010100001100",
   "01010111100000111011111001000010110001111110100001011001111111110100110010100001100",
   "01010111101100001100110011110101001100001101011010110111000110100001001000101001110",
   "01010111101100001100110011110101001100001101011010110111000110100001001000101001110",
   "01010111110111011110001110010111001010101110110001011101000000000000000100011100010",
   "01010111110111011110001110010111001010101110110001011101000000000000000100011100010",
   "01011000000010110000001000101011100000100100011110101111101001000101110110110111110",
   "01011000000010110000001000101011100000100100011110101111101001000101110110110111110",
   "01011000001110000010100010110101000001001000000111111010011010111001010011111000110",
   "01011000001110000010100010110101000001001000000111111010011010111001010011111000110",
   "01011000011001010101011100110110100000001011000001111011101010010100111111100001111",
   "01011000011001010101011100110110100000001011000001111011101010010100111111100001111",
   "01011000100100101000110110110010110001110110010101110001000010101011110101000000111",
   "01011000100100101000110110110010110001110110010101110001000010101011110101000000111",
   "01011000101111111100110000101100101010101011000100100100111011100000110001100111010",
   "01011000101111111100110000101100101010101011000100100100111011100000110001100111010",
   "01011000111011010001001010100110111111100010001011111100101010000001010010001010010",
   "01011000111011010001001010100110111111100010001011111100101010000001010010001010010",
   "01011001000110100110000100100100100101101100101010000111101110010010010110110100110",
   "01011001000110100110000100100100100101101100101010000111101110010010010110110100110",
   "01011001010001111011011110101000010010110011100010001111111100100000000101101010000",
   "01011001010001111011011110101000010010110011100010001111111100100000000101101010000",
   "01011001011101010001011000110100111100111000000000101010100010011111101001011011100",
   "01011001011101010001011000110100111100111000000000101010100010011111101001011011100",
   "01011001101000100111110011001101011010010011011111001010001001110011101111001001111",
   "01011001101000100111110011001101011010010011011111001010001001110011101111001001111",
   "01011001110011111110101101110100100001110111101001010001110110100011101001101100100",
   "01011001110011111110101101110100100001110111101001010001110110100011101001101100100",
   "01011001111111010110001000101101001010101110100000101001000011010101000111111001100",
   "01011001111111010110001000101101001010101110100000101001000011010101000111111001100",
   "01011010001010101110000011111010001100011010100001010000011010011001001110101011100",
   "01011010001010101110000011111010001100011010100001010000011010011001001110101011100",
   "01011010010110000110011111011110011110110110100101110111101100011100101101100100101",
   "01011010010110000110011111011110011110110110100101110111101100011100101101100100101",
   "01011010100001011111011011011100111010010110001100010100100101001100001001010111110",
   "01011010100001011111011011011100111010010110001100010100100101001100001001010111110",
   "01011010101100111000110111111000010111100101011001111010011101111100011101100011101",
   "01011010101100111000110111111000010111100101011001111010011101111100011101100011101",
   "01011010111000010010110100110011101111101000111111110011001110101000011010011011100",
   "01011010111000010010110100110011101111101000111111110011001110101000011010011011100",
   "01011011000011101101010010010001111011111110011111011000111101010011101010111101001",
   "01011011000011101101010010010001111011111110011111011000111101010011101010111101001",
   "01011011001111001000010000010101110110011100001110110000101100100100010010100111000",
   "01011011001111001000010000010101110110011100001110110000101100100100010010100111000",
   "01011011011010100011101111000010011001010001011101000110001001000011011000101111000",
   "01011011011010100011101111000010011001010001011101000110001001000011011000101111000",
   "01011011100101111111101110011010011111000110010111001000010110010101111100001000100",
   "01011011100101111111101110011010011111000110010111001000010110010101111100001000100",
   "01011011100101111111101110011010011111000110010111001000010110010101111100001000100",
   "01011011110001011100001110100001000010111100001011100111011011011110101110111110101",
   "01011011110001011100001110100001000010111100001011100111011011011110101110111110101",
   "01011011111100111001001111011001000000001101001111110011001111011010100000011011100",
   "01011011111100111001001111011001000000001101001111110011001111011010100000011011100",
   "01011100001000010110110001000101010010101101000011111011000101100111011110101010111",
   "01011100001000010110110001000101010010101101000011111011000101100111011110101010111",
   "01011100010011110100110011101000110110101000010111101110011011001001100001011111101",
   "01011100010011110100110011101000110110101000010111101110011011001001100001011111101",
   "01011100011111010011010111000110101000100101001110111110100100011100010010111111010",
   "01011100011111010011010111000110101000100101001110111110100100011100010010111111010",
   "01011100101010110010011011100001100101100011000110000001011100000100110001010000101",
   "01011100101010110010011011100001100101100011000110000001011100000100110001010000101",
   "01011100110110010010000000111100101010111010110110010101010010110011101001101101000",
   "01011100110110010010000000111100101010111010110110010101010010110011101001101101000",
   "01011101000001110010000111011010110110011110111011000101100001001010010011101110010",
   "01011101000001110010000111011010110110011110111011000101100001001010010011101110010",
   "01011101001101010010101110111111000110011011010101110000011010110011110110011100000",
   "01011101001101010010101110111111000110011011010101110000011010110011110110011100000",
   "01011101011000110011110111101100011001010101110010101110000100000100001010011011100",
   "01011101011000110011110111101100011001010101110010101110000100000100001010011011100",
   "01011101100100010101100001100101101110001101101101111000001001101110101110001011110",
   "01011101100100010101100001100101101110001101101101111000001001101110101110001011110",
   "01011101101111110111101100101110000100011100010111010010111011100111001001100001010",
   "01011101101111110111101100101110000100011100010111010010111011100111001001100001010",
   "01011101111011011010011001001000011011110100110111110111001001111101100010000000010",
   "01011101111011011010011001001000011011110100110111110111001001111101100010000000010",
   "01011110000110111101100110110111110100100100010101111101000110001000100111111011100",
   "01011110000110111101100110110111110100100100010101111101000110001000100111111011100",
   "01011110010010100001010101111111001111010001111010001000100110110000001001010011110",
   "01011110010010100001010101111111001111010001111010001000100110110000001001010011110",
   "01011110010010100001010101111111001111010001111010001000100110110000001001010011110",
   "01011110011110000101100110100001101100111110110011110110001111101001011101111110100",
   "01011110011110000101100110100001101100111110110011110110001111101001011101111110100",
   "01011110101001101010011000100010001111000110011110001001011101111001000101101111110",
   "01011110101001101010011000100010001111000110011110001001011101111001000101101111110",
   "01011110110101001111101100000011110111011110100100011011111000001011010111010111000",
   "01011110110101001111101100000011110111011110100100011011111000001011010111010111000",
   "01011111000000110101100001001001101000010111000111001101100011110111000100111000010",
   "01011111000000110101100001001001101000010111000111001101100011110111000100111000010",
   "01011111001100011011110111110110100100011010100000110110011110111100011111111101110",
   "01011111001100011011110111110110100100011010100000110110011110111100011111111101110",
   "01011111011000000010110000001101101110101101101010011000111111010011101110100000100",
   "01011111011000000010110000001101101110101101101010011000111111010011101110100000100",
   "01011111100011101010001010010010001010110000000000010101010111011101000101111111010",
   "01011111100011101010001010010010001010110000000000010101010111011101000101111111010",
   "01011111101111010010000110000110111100011011100111011110100001000110101001111011110",
   "01011111101111010010000110000110111100011011100111011110100001000110101001111011110",
   "01011111111010111010100011101111001000000101010001101111101101111001101111110110110",
   "01011111111010111010100011101111001000000101010001101111101101111001101111110110110",
   "01011111111010111010100011101111001000000101010001101111101101111001101111110110110",
   "01100000000110100011100011001101110010011100100011000011011110100011110001001011000",
   "01100000000110100011100011001101110010011100100011000011011110100011110001001011000",
   "01100000010010001101000100100110000000101011110110001011100000101101011001100110110",
   "01100000010010001101000100100110000000101011110110001011100000101101011001100110110",
   "01100000011101110111000111111010111000011000100001101001110011110011100110110010110",
   "01100000011101110111000111111010111000011000100001101001110011110011100110110010110",
   "01100000101001100001101101001111011111100010111100101010110101010101110011111010110",
   "01100000101001100001101101001111011111100010111100101010110101010101110011111010110",
   "01100000110101001100110100100110111100100110100100000000110100101100110010011011111",
   "01100000110101001100110100100110111100100110100100000000110100101100110010011011111",
   "01100001000000111000011110000100010110011001111111000000001110111101110111001000000",
   "01100001000000111000011110000100010110011001111111000000001110111101110111001000000",
   "01100001001100100100101001101010110100001111000100011101010010111110001001000100110",
   "01100001001100100100101001101010110100001111000100011101010010111110001001000100110",
   "01100001011000010001010111011101011101110010111111101010101101111001100110011001110",
   "01100001011000010001010111011101011101110010111111101010101101111001100110011001110",
   "01100001011000010001010111011101011101110010111111101010101101111001100110011001110",
   "01100001100011111110100111011111011011001110010101011001100000110001111000111100010",
   "01100001100011111110100111011111011011001110010101011001100000110001111000111100010",
   "01100001101111101100011001110011110101000101001000111001111111001000111011011011111",
   "01100001101111101100011001110011110101000101001000111001111111001000111011011011111",
   "01100001111011011010101110011101110100010111000000111101110111001011010110001111100",
   "01100001111011011010101110011101110100010111000000111101110111001011010110001111100",
   "01100010000111001001100101100000100010011111001100111011100011101111000001000000001",
   "01100010000111001001100101100000100010011111001100111011100011101111000001000000001",
   "01100010010010111000111110111111001001010100101001110010101000011001111101001001110",
   "01100010010010111000111110111111001001010100101001110010101000011001111101001001110",
   "01100010011110101000111010111100110011001010000111010001011000000110000011110010001",
   "01100010011110101000111010111100110011001010000111010001011000000110000011110010001",
   "01100010101010011001011001011100101010101110001100111011100110010110000111110101000",
   "01100010101010011001011001011100101010101110001100111011100110010110000111110101000",
   "01100010101010011001011001011100101010101110001100111011100110010110000111110101000",
   "01100010110110001010011010100001111011001011011111010010100011110000110100001100100",
   "01100010110110001010011010100001111011001011011111010010100011110000110100001100100",
   "01100011000001111011111110001111110000001000100100111110000101110110010100000110111",
   "01100011000001111011111110001111110000001000100100111110000101110110010100000110111",
   "01100011001101101110000100101001010101101000001011110110111010100101011010100101000",
   "01100011001101101110000100101001010101101000001011110110111010100101011010100101000",
   "01100011011001100000101101110001111000001001001110010010001000000101000100101010010",
   "01100011011001100000101101110001111000001001001110010010001000000101000100101010010",
   "01100011100101010011111001101100100100100110111000001101111000100111011000110111011",
   "01100011100101010011111001101100100100100110111000001101111000100111011000110111011",
   "01100011100101010011111001101100100100100110111000001101111000100111011000110111011",
   "01100011110001000111101000011100101000011000101100011111010011011011001100111100110",
   "01100011110001000111101000011100101000011000101100011111010011011011001100111100110",
   "01100011111100111011111010000101010001010010101010000001100010100001100010000101011",
   "01100011111100111011111010000101010001010010101010000001100010100001100010000101011",
   "01100100001000110000101110101001101101100101010001000110000101111100001110010100010",
   "01100100001000110000101110101001101101100101010001000110000101111100001110010100010",
   "01100100010100100110000110001101001011111101101000100110010100101011010001000110100",
   "01100100010100100110000110001101001011111101101000100110010100101011010001000110100",
   "01100100100000011100000000110010111011100101100011010110001011101110010111101010110",
   "01100100100000011100000000110010111011100101100011010110001011101110010111101010110",
   "01100100101100010010011110011110001100000011100101011000001011100000011100111111110",
   "01100100101100010010011110011110001100000011100101011000001011100000011100111111110",
   "01100100101100010010011110011110001100000011100101011000001011100000011100111111110",
   "01100100111000001001011111010010001101011011001001010010100100000010111000001000110",
   "01100100111000001001011111010010001101011011001001010010100100000010111000001000110",
   "01100101000100000001000011010010010000001100100101100101110000001110010010110000000",
   "01100101000100000001000011010010010000001100100101100101110000001110010010110000000",
   "01100101001111111001001010100001100101010101010010000100000000011111001000110101000",
   "01100101001111111001001010100001100101010101010010000100000000011111001000110101000",
   "01100101011011110001110101000011011110001111101101001010010101010011111001101101110",
   "01100101011011110001110101000011011110001111101101001010010101010011111001101101110",
   "01100101100111101011000010111011001100110011100001011010101001110011011001101111000",
   "01100101100111101011000010111011001100110011100001011010101001110011011001101111000",
   "01100101100111101011000010111011001100110011100001011010101001110011011001101111000",
   "01100101110011100100110100001100000011010101101010110111001110110001011010111111010",
   "01100101110011100100110100001100000011010101101010110111001110110001011010111111010",
   "01100101111111011111001000111001010100101000011100011111010110101000001011001001110",
   "01100101111111011111001000111001010100101000011100011111010110101000001011001001110",
   "01100110001011011010000001000110010011111011100101101101010010011101001011011011010",
   "01100110001011011010000001000110010011111011100101101101010010011101001011011011010",
   "01100110010111010101011100110110010100111100010111110101100000101000001111001001101",
   "01100110010111010101011100110110010100111100010111110101100000101000001111001001101",
   "01100110010111010101011100110110010100111100010111110101100000101000001111001001101",
   "01100110100011010001011100001100101011110101101011100111001101010011010101000011100",
   "01100110100011010001011100001100101011110101101011100111001101010011010101000011100",
   "01100110101111001101111111001100101101010000000110101110000101001010010110011101101",
   "01100110101111001101111111001100101101010000000110101110000101001010010110011101101",
   "01100110111011001011000101111001101110010010000001010101011010110001101111010111011",
   "01100110111011001011000101111001101110010010000001010101011010110001101111010111011",
   "01100111000111001000110000010111000100011111101011101100011110111011001001110010000",
   "01100111000111001000110000010111000100011111101011101100011110111011001001110010000",
   "01100111000111001000110000010111000100011111101011101100011110111011001001110010000",
   "01100111010011000110111110101000000101111011010011101100001100001111011110010111101",
   "01100111010011000110111110101000000101111011010011101100001100001111011110010111101",
   "01100111011111000101110000110000001001000101001010011110000110100101100011111101000",
   "01100111011111000101110000110000001001000101001010011110000110100101100011111101000",
   "01100111101011000101000110110010100100111011101010000100101110011101001111001110010",
   "10110110010100100011011111011010111010111110011100001111011101000100110000001110100",
   "10110110011010100011100000111010111100011110011101001011011101111001100100000101011",
   "10110110100000100011101011011011001111111111000011010000101011010000111001011101101",
   "10110110100000100011101011011011001111111111000011010000101011010000111001011101101",
   "10110110100110100011111110111100010000100010011100011000010000111101110110110001011",
   "10110110101100100100011011011110011001001100110000001110011011111000101000000010110",
   "10110110110010100101000001000010000101000100000000011101110101111000000011111100101",
   "10110110111000100101101111100111101111010000001000111011000011000001001100011110011",
   "10110110111110100110100111001111110010111010111111110000000000001100110111010111000",
   "10110111000100100111100111111010101011010000010101100111100011000011101010011011101",
   "10110111001010101000110001101000110011011101110101111000111011010000011000000010101",
   "10110111010000101010000100011010100110110011000110110011010101001001000111110001010",
   "10110111010000101010000100011010100110110011000110110011010101001001000111110001010",
   "10110111010110101011100000010000100000100001101001101001011101101111010111101011000",
   "10110111011100101101000101001010111011111100111010111101001000000111000010010011000",
   "10110111100010101110110011001010010100011010010010101010110100000100110101110100010",
   "10110111101000110000101010001111000101010001000100010101010110010100001000100100000",
   "10110111101110110010101010011001101001111010011111010001100001110100010111010110110",
   "10110111110100110100110011101010011101110001101110110001110010101110011010000001000",
   "10110111111010110111000110000001111100010011111010010001111010100001111010011111011",
   "10110111111010110111000110000001111100010011111010010001111010100001111010011111011",
   "10111000000000111001100001100000100001000000000101100010101101101010111011000001010",
   "10111000000110111100000110000110100111010111010000110101110010011111110111111001101",
   "10111000001100111110110011110100101010111100011001001001010001101000010001010010111",
   "10111000010011000001101010101011000111010100011000010011100111101100001001101101010",
   "10111000011001000100101010101010011000000110000101001111011000011100100101101010001",
   "10111000011111000111110011110010111000111010010100000111000011010101011001001111010",
   "10111000100101001011000110000101000101011011110110100000111001011000010000001000000",
   "10111000100101001011000110000101000101011011110110100000111001011000010000001000000",
   "10111000101011001110100001100001011001010111011011101010110100100001011100110100001",
   "10111000110001010010000110001000010000011011110000100110010000010110011011110000000",
   "10111000110111010101110011111010000110011001100000010100000100001110010111000110010",
   "10111000111101011001101010110111010111000011010100000000011110110100110111111110010",
   "10111001000011011101101011000000011110001101110011001111000011000111010001111011101",
   "10111001001001100001110100010101110111101111100100000110100110101100010101100100010",
   "10111001001111100110000110110111111111100001001011011101010001100110110111000101011",
   "10111001001111100110000110110111111111100001001011011101010001100110110111000101011",
   "10111001010101101010100010100111010001011101001101000100011111100011010101110101010",
   "10111001011011101111000111100100001001100000001011110101000010100000110001101001110",
   "10111001100001110011110101101111000011101000101001111011000110110100111011000111000",
   "10111001100111111000101101001000011011110111001001000010011000101100001011100101000",
   "10111001101101111101101101110000101110001110001010100010001011000101010010010000000",
   "10111001110100000010110111101000010110110010001111101001100000001001000011001010000",
   "10111001111010001000001010101111110001101001111001101011010010111110010101010100010",
   "10111001111010001000001010101111110001101001111001101011010010111110010101010100010",
   "10111010000000001101100111000111011010111101101010001010100010111010011101001010001",
   "10111010000110010011001100101111101110111000000011000110100000001110010000011011101",
   "10111010001100011000111011101001001001100101100111000110111010010000000000110010110",
   "10111010010010011110110011110100000111010100111001101000001111000010011010010111010",
   "10111010011000100100110101010001000100010110011111000111111100011000110011100000110",
   "10111010011110101011000000000000011100111100111101010000110010011000111011001110110",
   "10111010011110101011000000000000011100111100111101010000110010011000111011001110110",
   "10111010100100110001010100000010101101011100111011000111000111011010010011011011000",
   "10111010101010110111110001011000010010001101000001010101001101100011100100100010100",
   "10111010110000111110011000000001100111100101111010010111101001100101110111111100100",
   "10111010110111000101000111111111001010000010010010101001101011010110100110100011110",
   "10111010111101001100000001010001010101111110111000110001100111100111101001001010100",
   "10111011000011010011000011111000100111111010011101101101010011011110011000000010000",
   "10111011000011010011000011111000100111111010011101101101010011011110011000000010000",
   "10111011001001011010001111110101011100010101110100111110100001001001100111010110100",
   "10111011001111100001100101001000001111110011110100110111011110010110101110000111110",
   "10111011010101101001000011110001011110111001010110100111010100000110000101000111010",
   "10111011011011110000101011110001100110001101010110100110100111111111001011100110110",
   "10111011100001111000011101001001000010011000110100100011111111000100011111100110100",
   "10111011101000000000010111111000010000000110110011110000100010000111010111010001100",
   "10111011101000000000010111111000010000000110110011110000100010000111010111010001100",
   "10111011101110001000011011111111101100000100011011001100100011011100001001011010110",
   "10111011110100010000101001011111110011000000110101110100000110001110110010110001000",
   "10111011111010011001000000011001000001101101010010101011100111011000000101111101010",
   "10111100000000100001100000101011110100111101000101001100100111110011110100001001110",
   "10111100000110101010001010011000101001100101100101010010011000010111111100001000001",
   "10111100001100110010111101011111111100011110001111100110100111001101001101110111111",
   "10111100001100110010111101011111111100011110001111100110100111001101001101110111111",
   "10111100010010111011111010000010001010100000100101101110001110101001010000101101010",
   "10111100011001000100111111111111110000101000001110010110000101101010011001111001011",
   "10111100011111001110001111011001001011110010110101011111110001110101100001111001110",
   "10111100100101010111101000001110111001000000001100101110011010110110000110010111111",
   "10111100101011100001001010100001010101010010001011010011011111100000100110111111001",
   "10111100101011100001001010100001010101010010001011010011011111100000100110111111001",
   "10111100110001101010110110010000111101101100101110011011101100010111101011011001011",
   "10111100110111110100101011011110001111010101111001011011110011110100000000011101000",
   "10111100111101111110101010001001100111010101110101111101100111101111011011000000010",
   "10111101000100001000110010010011100010110110110100001100110100110011001110100010010",
   "10111101001010010011000011111100011111000101001011000011111111001010000110000010100",
   "10111101010000011101011111000100111001001111011000011001100000110101101101011101010",
   "10111101010000011101011111000100111001001111011000011001100000110101101101011101010",
   "10111101010110101000000011101101001110100110000001001100101001101000011010000110000",
   "10111101011100110010110001110101111100011011110001110010100000100011000000100001100",
   "10111101100010111101101001011111100000000101011110000011000110110111000110011000100",
   "10111101101001001000101010101010010110111010000001100110011100101101111110101011000",
   "10111101101111010011110101010110111110010010100000000001100111010100011111000100101",
   "10111101101111010011110101010110111110010010100000000001100111010100011111000100101",
   "10111101110101011111001001100101110011101010000101000011111000101011111100111010011",
   "10111101111011101010100111010111010100011110000100110011111001000000100000011010000",
   "10111110000001110110001110101011111110001101111011111100110001100100111100111000010",
   "10111110001000000001111111100100001110011011001111111011011001010100011100101011001",
   "10111110001110001101111010000000100010101001101111001011100010111010001111100000001",
   "10111110001110001101111010000000100010101001101111001011100010111010001111100000001",
   "10111110010100011001111110000001011000011111010001010101001100011111101010000100000",
   "10111110011010100110001011100111001101100011110111011001110001000000100101101111010",
   "10111110100000110010100010110010011111100001101100000001011011000110101111010000110",
   "10111110100110111111000011100011101100000101000011101000011001101011110011010010010",
   "10111110101101001011101101111011010000111100011100101100010110000010110111110000010",
   "10111110101101001011101101111011010000111100011100101100010110000010110111110000010",
   "10111110110011011000100001111001101011111000011111111001101011101001010001001011010",
   "10111110111001100101011111011111011010101100000000011001000001011111000010101101100",
   "10111110111111110010100110101100111011001011111011111100100101000111011000010000110",
   "10111111000101111111110111100010101011001111011011001101100111010001001001100110011",
   "10111111001100001101010010000001001000101111110001111001111010000111110101101111010",
   "10111111001100001101010010000001001000101111110001111001111010000111110101101111010",
   "10111111010010011010110110001000110001101000011111000001010001001101000101101110000",
   "10111111011000101000100011111010000011110111001101000011000010111011000110000011111",
   "10111111011110110110011011010101011101011011110010001011101011110000000110001001010",
   "10111111100101000100011100011011011100011000010000100010010011000011001100110111000",
   "10111111101011010010100111001100011110110000110110010110010001100010110001110110110",
   "10111111101011010010100111001100011110110000110110010110010001100010110001110110110",
   "10111111110001100000111011101001000010101011111110001100111001011100101010110100100",
   "10111111110111101111011001110001100110010010001111001111000000010000011100001100100",
   "10111111111101111110000001100110100111101110011101010110101010001011111100110110010",
   "11000000000100001100110011001000100101001101101001011100110111010010011100001100010",
   "11000000000100001100110011001000100101001101101001011100110111010010011100001100010",
   "11000000001010011011101110010111111100111111000001100111010010001110011010010101000",
   "11000000010000101010110011010101001101010100000001010110000000101110100001110101000",
   "11000000010110111010000010000000110100100000010001110001010101101101110010110001110",
   "11000000011101001001011010011011010000111001101001110111100101000111001110110011101",
   "11000000100011011000111100100101000000111000001110101010111001010101010101110011001",
   "11000000100011011000111100100101000000111000001110101010111001010101010101110011001",
   "11000000101001101000101000011110100010110110010011011111001010011101100011000101000",
   "11000000101111111000011110001000010101010000011010000111110111000111111010111000100",
   "11000000110110001000011101100010110110100101010011000101111111000011010111111110001",
   "11000000111100011000100110101110100101010101111101110101111111010110101001010010100",
   "11000001000010101000111001101100000000000101101000111101110000011110001111100110000",
   "11000001000010101000111001101100000000000101101000111101110000011110001111100110000",
   "11000001001000111001010110011011100101011001110010011010100101110111101011000101000",
   "11000001001111001001111100111101110011111010000111101111001111011010001000111101000",
   "11000001010101011010101101010011001010010000100110010001111100011101000001001001000",
   "11000001011011101011100111011100000111001001011011011010100000101100010100000110100",
   "11000001011011101011100111011100000111001001011011011010100000101100010100000110100",
   "11000001100001111100101011011001001001010011000100110000011010101011011001000010010",
   "11000001101000001101111001001010101111011110010000011000111100000110001100100101110",
   "11000001101110011111010000110001011000011101111101000101010011110001010000010111111",
   "11000001110100110000110010001101100011000111011010100000111001011000101011100000100",
   "11000001110100110000110010001101100011000111011010100000111001011000101011100000100",
   "11000001111011000010011101011111101110010010001001011111011010111110011100100110011",
   "11000010000001010100010010101000011000110111111100001011001100001000001101011101110",
   "11000010000111100110010001101000000001110100110110010011010110111100111001000011011",
   "11000010001101111000011010011111001000000111001101011010001110110010010100000000110",
   "11000010010100001010101101001110001010101111101001000011100100101011001000011011010",
   "11000010010100001010101101001110001010101111101001000011100100101011001000011011010",
   "11000010011010011101001001110101101000110001000011000010111101100101010101001111000",
   "11000010100000101111110000010110000001010000100111101010001010011001100001111110111",
   "11000010100111000010100000101111110011010101110101110111100001101011010111011111111",
   "11000010101101010101011011000011011110001010011111100100011011001011001110001100010",
   "11000010101101010101011011000011011110001010011111100100011011001011001110001100010",
   "11000010110011101000011111010001100000111010101001110011101101001001100010101110100",
   "11000010111001111011101101011010011010110100101101000000001011011100000001110100100",
   "11000011000000001111000101011110101011001001010101001011001000010100111011111110001",
   "11000011000110100010100111011110110001001011100010001010110111001100110010000010110",
   "11000011000110100010100111011110110001001011100010001010110111001100110010000010110",
   "11000011001100110110010011011011001100010000100111111001010000111110101011100010001",
   "11000011010011001010001001010100011011110000001110100010011010010111100111100011110",
   "11000011011001011110001001001010111111000100010010110011001011111000111001100000011",
   "11000011011111110010010010111111010101101001000110000111111011101110000010011010001",
   "11000011011111110010010010111111010101101001000110000111111011101110000010011010001",
   "11000011100110000110100110110001111110111101001110111011001001010110011000001011001",
   "11000011101100011011000100100011011010100001101000110100001011000010101011110000000",
   "11000011110010101111101100010100000111111001100100110101111101000110111111011101011",
   "11000011111001000100011110000100100110101010101001101101110011000000111110101101011",
   "11000011111001000100011110000100100110101010101001101101110011000000111110101101011",
   "11000011111111011001011001110101010110011100110100000010001010010011001000010111101",
   "11000100000101101110011111100110110110111010010110100001011111010100111101001000100",
   "11000100001100000011101111011001100111101111111010010001000011111000100011001111110",
   "11000100010010011001001001001110001000101100011110111011110111100101110001000001010",
   "11000100010010011001001001001110001000101100011110111011110111100101110001000001010",
   "11000100011000101110101101000100111001100001011011000001100010001011001111100100100",
   "11000100011111000100011010111110011010000010011100000101001111100101100111010111010",
   "11000100100101011010010010111011001010000101100110111100101101111101001000000001101",
   "11000100101011110000010100111011101001100011010111111111001101011001111101001001101",
   "11000100101011110000010100111011101001100011010111111111001101011001111101001001101",
   "11000100110010000110100001000000011000010110100011010100100001101111100001101001001",
   "11000100111000011100110111001001110110011100010101000100000101111111000011011001010",
   "11000100111110110011010111011000100011110100010001100100000001110001101000111111001",
   "11000101000101001010000001101101000000100000010101101000010000101010001011010000011",
   "11000101000101001010000001101101000000100000010101101000010000101010001011010000011",
   "11000101001011100000110110000111101100100100110110110001101011001111010100100011001",
   "11000101010001110111110100101001001000001000100011011101010010001101110111100101010",
   "11000101011000001110111101010001110011010100100011010011011011010011101111110101100",
   "11000101011110100110010000000010001110010100010111010111000000000011111101100000000",
   "11000101011110100110010000000010001110010100010111010111000000000011111101100000000",
   "11000101100100111101101100111010111001010101111010010100101110100011101110111111110",
   "11000101101011010101010011111100010100101001100000110010011100000001001010001010101",
   "11000101110001101101000101000111000000100001111001011110011001010011100111010011110",
   "11000101110001101101000101000111000000100001111001011110011001010011100111010011110",
   "11000101111000000101000000011011011101010100001101011110101001010110010000001100011",
   "11000101111110011101000101111010001011011000000000100000011001011100110101010111000",
   "11000110000100110101010101100011101011000111010001000111011011100011001011111100001",
   "11000110001011001101101111011000011100111110011000111101100010010111100110010111101",
   "11000110001011001101101111011000011100111110011000111101100010010111100110010111101",
   "11000110010001100110010011011001000001011100001101000001111111100000011010011001010",
   "11000110010111111111000001100101111001000001111101111001000011011101000110110001100",
   "11000110011110010111111001111111100100010011010111111011011111100011001011001101011",
   "11000110100100110000111100100110100011110110100011100110001001110111000101000001001",
   "11000110100100110000111100100110100011110110100011100110001001110111000101000001001",
   "11000110101011001010001001011011011000010100000101101001100011000001100011001010001",
   "11000110110001100011100000011110100010010110111111011001011110000001100100001111110",
   "11000110110111111101000001110000100010101100101110111100101001111011010001001111110",
   "11000110110111111101000001110000100010101100101110111100101001111011010001001111110",
   "11000110111110010110101101010001111010000101001111011100011101100100000111100111010",
   "11000111000100110000100011000011001001010010111001010100100101001100100101101000100",
   "11000111001011001010100011000100110001001010100010100010110010000111101011111000001",
   "11000111010001100100101101010111010010100011011110110110101100010000100110100101111",
   "11000111010001100100101101010111010010100011011110110110101100010000100110100101111",
   "11000111010111111111000001111011001110010111100000000001100101101110110010000011010",
   "11000111011110011001100000110001000101100010110110000110010000011000101100110101001",
   "11000111100100110100001001111001011001000100001111101000110101010101101011000011101",
   "11000111100100110100001001111001011001000100001111101000110101010101101011000011101",
   "11000111101011001110111101010100101001111100111001111110101110011110111101110001110",
   "11000111110001101001111011000011011001010000100001011110100010000000100001100100100",
   "11000111111000000101000011000110001000000101010001101111111111111001100111101000101",
   "11000111111110100000010101011101010111100011110101111100000001011101101100100111010",
   "11000111111110100000010101011101010111100011110101111100000001011101101100100111010",
   "11001000000100111011110010001001101000110111011000111100101010110101110000011110010",
   "11001000001011010111011001001011011101001101100101101101001110100010100010110100010",
   "11001000010001110011001010100011010101110110100111011010010010111111110111000010101",
   "11001000010001110011001010100011010101110110100111011010010010111111110111000010101",
   "11001000011000001111000110010001110100000101001001110001111010001001010011110101100",
   "11001000011110101011001100010111011001001110011001010011101011000000110001100011000",
   "11001000100101000111011100110100100110101010000011100000111101010110111010111110000",
   "11001000100101000111011100110100100110101010000011100000111101010110111010111110000",
   "11001000101011100011110111101001111101110010010111001101000111010110000100010001011",
   "11001000110010000000011100111000000000000100000100101101101101001111101011101010101",
   "11001000111000011101001100011111001110111110011110001010110011001100110111101000100",
   "11001000111110111010000110100000001100000011010111101111010001000010000110011110010",
   "11001000111110111010000110100000001100000011010111101111010001000010000110011110010",
   "11001001000101010111001010111011011000110111000111111001001000000110100011000011111",
   "11001001001011110100011001110001010111000000100111101001111011001111010010101100010",
   "11001001010010010001110011000010101000001001010010110111001000101110110000000001001",
   "11001001010010010001110011000010101000001001010010110111001000101110110000000001001",
   "11001001011000101111010110101111101101111101001000011010100110011000100111000011110",
   "11001001011111001101000100111001001010001010101010100010111111101010100110011010000",
   "11001001100101101010111101011111011110100010111111000100010101111010011001101101110",
   "11001001100101101010111101011111011110100010111111000100010101111010011001101101110",
   "11001001101100001001000000100011001100111001101111101000100010101001000001101101000",
   "11001001110010100111001110000100110111000101001001111111111011111011111101111000100",
   "11001001111001000101100110000100111110111110000000010001111010111100011100010101010",
   "11001001111111100100001000100100000110011111101001001101100100011101000011110111010",
   "11001001111111100100001000100100000110011111101001001101100100011101000011110111010",
   "11001010000110000010110101100010101111101000000000011010010011100110001100111111110",
   "11001010001100100001101101000001011100010111100110101000100110101001011110001110011",
   "11001010010011000000101111000000101110110001100010000010101101111100100000000100000",
   "11001010010011000000101111000000101110110001100010000010101101111100100000000100000",
   "11001010011001011111111011100001001000111011011110011101011100111011011101100000000",
   "11001010011111111111010010100011001100111101101101101000111101010011100101011111000",
   "11001010100110011110110100000111011101000011000111100001100100010110000010000111100",
   "11001010100110011110110100000111011101000011000111100001100100010110000010000111100",
   "11001010101100111110100000001110011011011001001010100000101010010011011010010101001",
   "11001010110011011110010110111000101010001111111011101101100100000000010010111000010",
   "11001010111001111110011000000110101011111010000111001110011110100011000011011110010",
   "11001010111001111110011000000110101011111010000111001110011110100011000011011110010",
   "11001011000000011110100011111001000010101101000000011001011101001011010101000000100",
   "11001011000110111110111010010000010001000000100010000101011001010011011101111000001",
   "11001011001101011111011011001100111001001111001110111011000100101100010001011010100",
   "11001011001101011111011011001100111001001111001110111011000100101100010001011010100",
   "11001011010100000000000110101111011101110110010001100110001101110011010111100010011",
   "11001011011010100000111100111000100001010101011101000110100110010100100001110100100",
   "11001011100001000001111101101000100110001111001101000001001011110110010011001000111",
   "11001011100001000001111101101000100110001111001101000001001011110110010011001000111",
   "11001011100111100011001001000000001111001000100101110001010010110010001111001110011",
   "11001011101110000100011110111111111110101001010100111001110011011001000111011100101",
   "11001011110100100101111111101000010111011011110001010110011001000011011010001110010",
   "11001011110100100101111111101000010111011011110001010110011001000011011010001110010",
   "11001011111011000111101010111001111100001100111011101100110011101110011010100000100",
   "11001100000001101001100000110101001111101100011110011110001011100110010100111010000",
   "11001100001000001011100001011010110100101100101110011000010110111101100111111100111",
   "11001100001000001011100001011010110100101100101110011000010110111101100111111100111",
   "11001100001110101101101100101011001110000010101010100111010010010010000101001101100",
   "11001100010101010000000010100110111110100101111101000110011010011111110000111011011",
   "11001100011011110010100011001110101001010000111010110010001001100010010101111011000",
   "11001100011011110010100011001110101001010000111010110010001001100010010101111011000",
   "11001100100010010101001110100010110001000000100011111001010101000101000011100111000",
   "11001100101000111000000100100011111000110100100100001110101111100001101100000000100",
   "11001100101111011011000101010010100011101111010011011010101011001110110111101001101",
   "11001100101111011011000101010010100011101111010011011010101011001110110111101001101",
   "11001100110101111110010000101111010100110101110101001100011111111110000101011100101",
   "11001100111100100001100110111010101111001111111001101100010010101001101100100010110",
   "11001101000011000101000111110101010110000111111101101100011111010011010110010010100",
   "11001101000011000101000111110101010110000111111101101100011111010011010110010010100",
   "11001101001001101000110011011111101100101011001010111011100101010011000110100010011",
   "11001101010000001100101001111010010110001001011000010101110101110111101000100000000",
   "11001101010110110000101011000101110101110101001010010111000100110111110110011111001",
   "11001101010110110000101011000101110101110101001010010111000100110111110110011111001",
   "11001101011101010100110111000010101111000011110011001100011011110110010010111001010",
   "11001101100011111001001101110001100101001101010011000110001111010110101000111010010",
   "11001101101010011101101111010010111011101100011000101001110110100101101011011000111",
   "11001101101010011101101111010010111011101100011000101001110110100101101011011000111",
   "11001101110001000010011011100111010101111110100001000011100101010100001000100001000",
   "11001101110111100111010010101111010111100011111000011000101000000100101000110110110",
   "11001101111110001100010100101011100011111111011001111001000010101101010000011111001",
   "11001101111110001100010100101011100011111111011001111001000010101101010000011111001",
   "11001110000100110001100001011100011110110110110000010001110001001100111000111110101",
   "11001110001011010110111001000010101011110010010101111110101010110100111011000010100",
   "11001110010001111100011011011110101110011101010101011100100111100111011110101101011",
   "11001110010001111100011011011110101110011101010101011100100111100111011110101101011",
   "11001110011000100010001000110001001010100101101001011011101000001010101001000010101",
   "11001110011111001000000000111010100011111011111101010000111111110000111110010100001",
   "11001110011111001000000000111010100011111011111101010000111111110000111110010100001",
   "11001110100101101110000011111011011110010011101101001001100000110111101111110100100",
   "11001110101100010100010001110100011101100011000110011011101011111011001100011001010",
   "11001110110010111010101010100110000101100011000111111010000000100001001010111000010",
   "11001110110010111010101010100110000101100011000111111010000000100001001010111000010",
   "11001110111001100001001110010000111010001111100010000101010000111010100101110100110",
   "11001111000000000111111100110101011111100110110111011110110111111011111111101110000",
   "11001111000110101110110110010100011001101010011100111011010001001101100111001101110",
   "11001111000110101110110110010100011001101010011100111011010001001101100111001101110",
   "11001111001101010101111010101110001100011110011001110100010011110011010010110001011",
   "11001111010011111101001010000011011100001001101000011011101111001100101011010001010",
   "11001111011010100100100100010100101100110101110110001101101010101101111101001110001",
   "11001111011010100100100100010100101100110101110110001101101010101101111101001110001",
   "11001111100001001100001001100010100010101111100100000011000111010001101000001110011",
   "11001111100111110011111001101101100010000110000110100100100011100011100100011001100",
   "11001111100111110011111001101101100010000110000110100100100011100011100100011001100",
   "11001111101110011011110100110110001111001011100110011100100010100101110101101000110",
   "11001111110101000011111010111101001110010101000000101010010100101111100100100000001",
   "11001111111011101100001100000011000011111010000110110100100011000110010100110000100",
   "11001111111011101100001100000011000011111010000110110100100011000110010100110000100",
   "11010000000010010100101000001000010100010101011111011011111101010010010001100000101",
   "11010000001000111101001111001101100100000100100110001110001001101101100111000001110",
   "11010000001111100110000001010011010111100111101100011000011000001111100010011100010",
   "11010000001111100110000001010011010111100111101100011000011000001111100010011100010",
   "11010000010110001110111110011010010011100001111000111010010111010011001111011101010",
   "11010000011100111000000110100010111100011001001000111001001011011011001100011011111",
   "11010000011100111000000110100010111100011001001000111001001011011011001100011011111",
   "11010000100011100001011001101101110110110110001111110010001001010001001101001001110",
   "11010000101010001010110111111011100111100100110111101101110010000011100100101001101",
   "11010000110000110100100001001100110011010011100001110010110010011111101110101110100",
   "11010000110000110100100001001100110011010011100001110010110010011111101110101110100",
   "11010000110111011110010101100001111110110011100110011001000100001010110001100010010",
   "11010000111110001000010100111011101110111001010101011100110001011000010000000000101",
   "11010000111110001000010100111011101110111001010101011100110001011000010000000000101",
   "11010001000100110010011111011010101000011011110110110001011011011111100101110000110",
   "11010001001011011100110100111111010000010101001010010101000011110000100101001110101",
   "11010001010010000111010101101010001011100010001000100011010110100111010000111011011",
   "11010001010010000111010101101010001011100010001000100011010110100111010000111011011",
   "11010001011000110010000001011011111111000010100010101000111001011111101000101101101",
   "11010001011111011100111000010101001111111001000010110110011011001001100100000001100",
   "11010001100110000111111010010110100011001011001100110100000110011101010010001011010",
   "11010001100110000111111010010110100011001011001100110100000110011101010010001011010",
   "11010001101100110011000111100000011110000001011101110100110111110000111001110100010",
   "11010001110011011110011111110011100101100111001101001001110100101111010000101111100",
   "11010001110011011110011111110011100101100111001101001001110100101111010000101111100",
   "11010001111010001010000011010000011111001010101100010101100110110000100101010110101",
   "11010010000000110101110001110111101111111101000111011111110111110101010011000101011",
   "11010010000111100001101011101001111101010010100101101000110010000011011011001100100",
   "11010010000111100001101011101001111101010010100101101000110010000011011011001100100",
   "11010010001110001101110000100111101100100010001000111100100001100110111011011110000",
   "11010010010100111010000000110001100011000101101111000110111001010101011100010011010",
   "11010010010100111010000000110001100011000101101111000110111001010101011100010011010",
   "11010010011011100110011100001000000110011010010001100110111001110101101111111000000",
   "11010010100010010011000010101011111011111111100110000010011011001011011100000101100",
   "11010010101000111111110100011101101001011000011110011001111001000111001001000001000",
   "11010010101000111111110100011101101001011000011110011001111001000111001001000001000",
   "11010010101111101100110001011101110100001010101001011100000001111011101101110010111",
   "11010010110110011001111001101101000001111110110010111001100111111000110101110011000",
   "11010010110110011001111001101101000001111110110010111001100111111000110101110011000",
   "11010010111101000111001101001011111000100000100011111001010101001011011000001000001",
   "11010011000011110100101011111010111101011110100011001011100010100011111011100010110",
   "11010011001010100010010101111010110110101010010101011110010000100100000000111001010",
   "11010011001010100010010101111010110110101010010101011110010000100100000000111001010",
   "11010011010001010000001011001100001001111000011101110001000011010010001110010101011",
   "11010011010111111110001011101111011101000000011101101001000000110101110101100111100",
   "11010011010111111110001011101111011101000000011101101001000000110101110101100111100",
   "11010011011110101100010111100101010101111100110101100100110010011010001111110100101",
   "11010011100101011010101110101110011010101011000101010000100111111010101000111111010",
   "11010011100101011010101110101110011010101011000101010000100111111010101000111111010",
   "11010011101100001001010001001011010001001011101011111010011110010110010110001010111",
   "11010011110010110111111110111100011111100010001000100110001000101110010000100000110",
   "11010011111001100110111000000010101011110100111010100001011011101011110000000010110",
   "11010011111001100110111000000010101011110100111010100001011011101011110000000010110",
   "11010100000000010101111100011110011100001101100001011000011011110001100000111011111",
   "11010100000111000101001100010000010110111000011101101001101110010110101110000011011",
   "11010100000111000101001100010000010110111000011101101001101110010110101110000011011",
   "11010100001101110100100111011001000010000101010000111010101101001100111011101101101",
   "11010100010100100100001101111001000100000110011110001011111100110001001101101010010",
   "11010100011011010011111111110001000011010001101010001101100101001000110011010010010",
   "11010100011011010011111111110001000011010001101010001101100101001000110011010010010",
   "11010100100010000011111101000001100101111111011011110011101101101001110101010001010",
   "11010100101000110100000101101011010010101011011100001010111011010000011111110110101",
   "11010100101000110100000101101011010010101011011100001010111011010000011111110110101",
   "11010100101111100100011001101110101111110100010111001100110001100001000101000011011",
   "11010100110110010100111001001100100011111011111011110100010110010111010010001010101",
   "11010100110110010100111001001100100011111011111011110100010110010111010010001010101",
   "11010100111101000101100100000101010101100110111100010010111000100011010100000101100",
   "11010101000011110110011010011001101011011101001110100100011000110101000101111001010",
   "11010101001010100111011100001010001100001001101100100100010101110110000101011011000",
   "11010101001010100111011100001010001100001001101100100100010101110110000101011011000",
   "11010101010001011000101001010111011110011010010100100010011010110010001001011001110",
   "11010101011000001010000010000010001001000000001001010111010000101111110101000011111",
   "11010101011000001010000010000010001001000000001001010111010000101111110101000011111",
   "11010101011110111011100110001010110010101111010010111001010010111000100100111101010",
   "11010101100101101101010101110010000010011110111110010001100101010001010001000011000",
   "11010101100101101101010101110010000010011110111110010001100101010001010001000011000",
   "11010101101100011111010000111000011111001001011110010000101110100011011111111100010",
   "11010101110011010001010111011110101111101100001011100011110100011000000111100010110",
   "11010101111010000011101001100101011011000111100101001001011010100011010111001001001",
   "11010101111010000011101001100101011011000111100101001001011010100011010111001001001",
   "11010110000000110110000111001101001000011111010000100110100101000011000111010100101",
   "11010110000111101000110000010110011110111001111010011011111100101111101011111110110",
   "11010110000111101000110000010110011110111001111010011011111100101111101011111110110",
   "11010110001110011011100101000010000101100001010110011010110110111111100100111001000",
   "11010110010101001110100101010000100011100010011111111010011111111110101001010110101",
   "11010110010101001110100101010000100011100010011111111010011111111110101001010110101",
   "11010110011100000001110001000010100000001101011010001101000111111001001011011110000",
   "11010110100010110101001000011000100010110101010000110101010010111011001111110010001",
   "11010110100010110101001000011000100010110101010000110101010010111011001111110010001",
   "11010110101001101000101011010011010010110000010111111011001100000100110110000000001",
   "11010110110000011100011001110011010111011000001100100001111010110011001111101010101",
   "11010110110111010000010011111001011000001001010100111100111011100000000001101011110",
   "11010110110111010000010011111001011000001001010100111100111011100000000001101011110",
   "11010110111110000100011001100101111100100011100001000101011010110110001101110000001",
   "11010111000100111000101010111001101100001001101010101111110011111110000000110000011",
   "11010111000100111000101010111001101100001001101010101111110011111110000000110000011",
   "11010111001011101101000111110101001110100001110110000001010001011111100011010101000",
   "11010111010010100001110000011001001011010101010001100101010001011101001001110110011",
   "11010111010010100001110000011001001011010101010001100101010001011101001001110110011",
   "11010111011001010110100100100110001010010000010111000011001100000101100001001101011",
   "11010111100000001011100100011100110011000010101011010011111101011110010101110011100",
   "11010111100000001011100100011100110011000010101011010011111101011110010101110011100",
   "11010111100111000000101111111101101101011110111110110111110010000111110010010010000",
   "11010111101101110110000111001001100001011011001110001011110110011001010011100111001",
   "11010111101101110110000111001001100001011011001110001011110110011001010011100111001",
   "11010111110100101011101010000000110110110000100010000000001000111000010000001111110",
   "11010111111011100001011000100100010101011011001111101101001111101000110000000101100",
   "11010111111011100001011000100100010101011011001111101101001111101000110000000101100",
   "11011000000010010111010010110100100101011010111001101010010000011001010011001010100",
   "11011000001001001101011000110010001110110010001111100010101011101001100100111110101",
   "11011000010000000011101010011101111001100111001110101100011010101100111010100011101",
   "11011000010000000011101010011101111001100111001110101100011010101100111010100011101",
   "11011000010110111010000111111000001110000011000010011101110000101000111001010101110",
   "11011000011101110000110001000001110100010010000100100011011110010000100101001001000",
   "11011000011101110000110001000001110100010010000100100011011110010000100101001001000",
   "11011000100100100111100101111011010100100011111101010110111000111100110011011101111",
   "11011000101011011110100110100101010111001011100100010100000100100010000010101000101",
   "11011000101011011110100110100101010111001011100100010100000100100010000010101000101",
   "11011000110010010101110011000000100100011111000000010000000000000100010011000111111",
   "11011000111001001101001011001101100100110111100111101110110101101001100001110001100",
   "11011000111001001101001011001101100100110111100111101110110101101001100001110001100",
   "11011001000000000100101111001101000000110010000001011010001101001011000001100000100",
   "11011001000110111100011110111111100000101110000100010111100010000110010011010010100",
   "11011001000110111100011110111111100000101110000100010111100010000110010011010010100",
   "11011001001101110100011010100101101101001110111000011110011100001101111011001101001",
   "11011001010100101100100010000000001110111010110110101111001011011010110001100110111",
   "11011001010100101100100010000000001110111010110110101111001011011010110001100110111",
   "11011001011011100100110101001111101110011011101001101001000110011110001111010100001",
   "11011001100010011101010100010100110100011110001101100001001100110101110100000001100",
   "11011001100010011101010100010100110100011110001101100001001100110101110100000001100",
   "11011001101001010101111111010000001001110010110000111000101011100000100110001000100",
   "11011001110000001110110110000010010111001100110100110011100100110111001011010001110",
   "11011001110000001110110110000010010111001100110100110011100100110111001011010001110",
   "11011001110111000111111000101100000101100011001101001111011011100110011000111110101",
   "11011001111110000001000111001101111101110000000001011010000000101101011100111001000",
   "11011001111110000001000111001101111101110000000001011010000000101101011100111001000",
   "11011010000100111010100001101000101000110000101100001000000100011111111100001110111",
   "11011010001011110100000111111100101111100101111100001100001010101100001010000100111",
   "11011010001011110100000111111100101111100101111100001100001010101100001010000100111",
   "11011010010010101101111010001010111011010011110100101101100001100110010100010000001",
   "11011010011001100111111000010011110101000001101101011110111100011001000110110000000",
   "11011010011001100111111000010011110101000001101101011110111100011001000110110000000",
   "11011010100000100010000010011000000101111010010011010101110000011100000101100011010",
   "11011010100111011100011000011000010111001011101000100000110101110000011100111101011",
   "11011010101110010110111010010101010010000111000100111111101010100100101000100100101",
   "11011010101110010110111010010101010010000111000100111111101010100100101000100100101",
   "11011010110101010001101000001111100000000001010110111001011001111111010001000111001",
   "11011010111100001100100010000111101010010010100010110100000101110010000001011110100",
   "11011010111100001100100010000111101010010010100010110100000101110010000001011110100",
   "11011011000011000111100111111110011010010110000100001011110011010100110011011100110",
   "11011011001010000010111001110100011001101010101101101001111011101001110100100010010",
   "11011011001010000010111001110100011001101010101101101001111011101001110100100010010",
   "11011011010000111110010111101010010001110010101001011100011110101011000011101000101",
   "11011011010111111010000001100000101100010011011001101101011001100001101000001100111",
   "11011011010111111010000001100000101100010011011001101101011001100001101000001100111",
   "11011011011110110101110111011000010010110101111000111010000000000111100011101110101",
   "11011011100101110001111001010001101111000110011010001010011001110100011110011111001",
   "11011011100101110001111001010001101111000110011010001010011001110100011110011111001",
   "11011011101100101110000111001101101010110100101001101001000001010101110000100000100",
   "11011011101100101110000111001101101010110100101001101001000001010101110000100000100",
   "11011011110011101010100001001100101111110011101100111010000111110010100111111011100",
   "11011011111010100111000111001111100111111010000011010011011010111100101101111010110",
   "11011011111010100111000111001111100111111010000011010011011010111100101101111010110",
   "11011100000001100011111001010110111101000001100110010011101110101101101011011101000",
   "11011100001000100000110111100011011001000111101001111010101001110010001111011010001",
   "11011100001000100000110111100011011001000111101001111010101001110010001111011010001",
   "11011100001111011110000001110101100110001100111101000000010101100011010111011010010",
   "11011100010110011011011000001110001110010101101001101101010001001101111101000101000",
   "11011100010110011011011000001110001110010101101001101101010001001101111101000101000",
   "11011100011101011000111010101101111011101001010101110010001000001001101001011000011",
   "11011100100100010110101001010101011000010011000010111111101011011111001111110111010",
   "11011100100100010110101001010101011000010011000010111111101011011111001111110111010",
   "11011100101011010100100100000101001110100001001111011110101110111111010011101100011",
   "11011100110010010010101010111110001000100101110110001000001001001001011000100001010",
   "11011100110010010010101010111110001000100101110110001000001001001001011000100001010",
   "11011100111001010000111110000000110000110110001110111100110110100100100001001110101",
   "11011101000000001111011101001101110001101011001111011110000000101001011110110110001",
   "11011101000000001111011101001101110001101011001111011110000000101001011110110110001",
   "11011101000111001110001000100101110101100001001011000101000111011111010001110110101",
   "11011101001110001101000000001001100110110111110011011100001111001010100000010111110",
   "11011101001110001101000000001001100110110111110011011100001111001010100000010111110",
   "11011101010101001100000011111001110000010010011000110110010000010000000011101101000",
   "11011101011100001011010011110110111100010111101010100111001011101011101111110110000",
   "11011101011100001011010011110110111100010111101010100111001011101011101111110110000",
   "11011101100011001010110000000001110101110001110111011100100001111011010111101110110",
   "11011101101010001010011000011011000111001110101101110101101101011110110000111111011",
   "11011101101010001010011000011011000111001110101101110101101101011110110000111111011",
   "11011101110001001010001101000011011011011111011100011100100000101101011010001010110",
   "11011101111000001010001101111011011101011000110010011101100111000010000110011100110",
   "11011101111000001010001101111011011101011000110010011101100111000010000110011100110",
   "11011101111111001010011011000011110111110011000000000001001001011101010010000001011",
   "11011110000110001010110100011101010101101001110110100011010110011110100010010011111",
   "11011110000110001010110100011101010101101001110110100011010110011110100010010011111",
   "11011110001101001011011010001000100001111100101001001101001101010101110101011101000",
   "11011110001101001011011010001000100001111100101001001101001101010101110101011101000",
   "11011110010100001100001100000110000111101110001101001101001100101101000100011101000",
   "11011110011011001101001010010110110010000100111010010000000100101010011011100110101",
   "11011110011011001101001010010110110010000100111010010000000100101010011011100110101",
   "11011110100010001110010100111011001100001010101010111001101100001100001100110011000",
   "11011110101001001111101011110100000001001100111100111101111001111110011111100100010",
   "11011110101001001111101011110100000001001100111100111101111001111110011111100100010",
   "11011110110000010001001111000001111100011100110001111001100000101011100010101011111",
   "11011110110111010010111110100101101001001110101111001011001110100111000011010101101",
   "11011110110111010010111110100101101001001110101111001011001110100111000011010101101",
   "11011110111110010100111010011111110010111010111110101100110000110101001101111101110",
   "11011111000101010111000010110001000100111101001111001011111001101101111100111111010",
   "11011111000101010111000010110001000100111101001111001011111001101101111100111111010",
   "11011111001100011001010111011010001010110100110100100011101010111100111001101110000",
   "11011111010011011011111000011011110000000100101000010101100010111110110011111001110",
   "11011111010011011011111000011011110000000100101000010101100010111110110011111001110",
   "11011111011010011110100101110110100000010011001010000010101101111100110100011001101",
   "11011111011010011110100101110110100000010011001010000010101101111100110100011001101",
   "11011111100001100001011111101011000111001010011111100101011010000110001111101011101",
   "11011111101000100100100101111010010000011000010101101010001111101001011100111000000",
   "11011111101000100100100101111010010000011000010101101010001111101001011100111000000",
   "11011111101111100111111000100100100111101110000000001001101100001100010110001111010",
   "11011111110110101011010111101010111001000000011010100001100001100101001000000001100",
   "11011111110110101011010111101010111001000000011010100001100001100101001000000001100",
   "11011111111101101111000011001101110000001000001000001110011000010011110010110110000",
   "11100000000100110010111011001101111001000001010101000101010101011101000110101110011",
   "11100000000100110010111011001101111001000001010101000101010101011101000110101110011",
   "11100000001011110110111111101011111111101011110101101101100100000111011100001010001",
   "11100000010010111011010000101000110000001011000111111010000010011010010000100101011",
   "11100000010010111011010000101000110000001011000111111010000010011010010000100101011",
   "11100000011001111111101110000100110110100110010011000011010010000000101011110110101",
   "11100000011001111111101110000100110110100110010011000011010010000000101011110110101",
   "11100000100001000100011000000000111111001000001000100001001100001111110100010011000",
   "11100000101000001001001110011101110101111111000100000100111001110001010111001100010",
   "11100000101000001001001110011101110101111111000100000100111001110001010111001100010",
   "11100000101111001110010001011100000111011101001100010010101101110011001011011111011",
   "11100000110110010011100000111100011111111000010010111100000100111100010100110100101",
   "11100000110110010011100000111100011111111000010010111100000100111100010100110100101",
   "11100000111101011000111100111111101011101001110101011001100111101000001100110110100",
   "11100001000100011110100101100110010111001110111101000101010000001000011001010000010",
   "11100001000100011110100101100110010111001110111101000101010000001000011001010000010",
   "11100001001011100100011010110001001111001000011111110100010100001101110100100111010",
   "11100001001011100100011010110001001111001000011111110100010100001101110100100111010",
   "11100001010010101010011100100000111111111011000000010001110010011001110000101111001",
   "11100001011001110000101010110110010110001110101110011000100010110111011000111011000",
   "11100001011001110000101010110110010110001110101110011000100010110111011000111011000",
   "11100001100000110111000101110001111110101111100111101101101011111110011010111001101",
   "11100001100111111101101101010100100110001101010111111010111010011111011101010000000",
   "11100001100111111101101101010100100110001101010111111010111010011111011101010000000",
   "11100001101111000100100001011110111001011011011001001000111101011010101010001100101",
   "11100001110110001011100010010001100101010000110100011010000101100001010101111000000",
   "11100001110110001011100010010001100101010000110100011010000101100001010101111000000",
   "11100001111101010010101111101101010110101000100010000100101000100011000111001011000",
   "11100001111101010010101111101101010110101000100010000100101000100011000111001011000",
   "11100010000100011010001001110010111010100001001010001101101000000111001010011111000",
   "11100010001011100001110000100010111101111101000101000011011100010010010101101111110",
   "11100010001011100001110000100010111101111101000101000011011100010010010101101111110",
   "11100010010010101001100011111110001110000010011011011000100001111010100101010001111",
   "11100010011001110001100100000101010111111011000110111110001100101000011001000101111",
   "11100010011001110001100100000101010111111011000110111110001100101000011001000101111",
   "11100010100000111001110000111001001000110100110010111111011100100110111010011001010",
   "11100010101000000010001010011010001110000000111100011011111000000011010001001110010",
   "11100010101000000010001010011010001110000000111100011011111000000011010001001110010",
   "11100010101111001010110000101001010100110100110010100010101000011011110010001001101",
   "11100010101111001010110000101001010100110100110010100010101000011011110010001001101",
   "11100010110110010011100011100111001010101001010111001101011011011111101100010000111",
   "11100010111101011100100011010100011100111011011111011011100111111111111111100101011",
   "11100010111101011100100011010100011100111011011111011011100111111111111111100101011",
   "11100011000100100101101111110001111001001011110011101101010110010010000100010111111",
   "11100011001011101111001001000000001100111110110000011110101100100100101011110010001",
   "11100011001011101111001001000000001100111110110000011110101100100100101011110010001",
   "11100011010010111000101111000000000101111100100110100010111111001000000010011110100",
   "11100011010010111000101111000000000101111100100110100010111111001000000010011110100",
   "11100011011010000010100001110010010001110001011011100000000100001001011101111101001",
   "11100011100001001100100001010111011110001101001010001001101011100011011101011111100",
   "11100011100001001100100001010111011110001101001010001001101011100011011101011111100",
   "11100011101000010110101101110000011001000011100010111100111010100010100111101000000",
   "11100011101111100001000110111101110000001100001100011011101011000000001101010110100",
   "11100011101111100001000110111101110000001100001100011011101011000000001101010110100",
   "11100011110110101011101101000000010001100010100011101000001110110010111100010000110",
   "11100011110110101011101101000000010001100010100011101000001110110010111100010000110",
   "11100011111101110110011111111000101011000101111100100000110110110110101000111111100",
   "11100100000101000001011111100111101010111001100010011011011110001011011011011111001",
   "11100100000101000001011111100111101010111001100010011011011110001011011011011111001",
   "11100100001100001100101100001101111111000100011000100001011000101101000110101011110",
   "11100100010011011000000101101100010101110001011010001011000110000011010101011001111",
   "11100100010011011000000101101100010101110001011010001011000110000011010101011001111",
   "11100100011010100011101100000011011101001111011011011100001000001011010110010011011",
   "11100100011010100011101100000011011101001111011011011100001000001011010110010011011",
   "11100100100001101111011111010100000011110001001001011110111101111011110000111001100",
   "11100100101000111011011111011110110111101101001011000001000001100011001101110100011",
   "11100100101000111011011111011110110111101101001011000001000001100011001101110100011",
   "11100100110000000111101100100100100111011110000000101110101011000010011100100010000",
   "11100100110000000111101100100100100111011110000000101110101011000010011100100010000",
   "11100100110111010100000110100110000001100010000101101111010110100010100000111101100",
   "11100100111110100000101101100011110100011011110000000001101110100111110011100001000",
   "11100100111110100000101101100011110100011011110000000001101110100111110011100001000",
   "11100101000101101101100001011110101110110001010000110111111010100010011110001011000",
   "11100101001100111010100010010111011111001100110101010011110000011101000001011100000",
   "11100101001100111010100010010111011111001100110101010011110000011101000001011100000",
   "11100101010100000111110000001110110100011100100110100011001011101001101100000101011",
   "11100101010100000111110000001110110100011100100110100011001011101001101100000101011",
   "11100101011011010101001011000101011101010010101010011100100110101111010000101101111",
   "11100101100010100010110010111100001000100101000011111011011001110110000100010111101",
   "11100101100010100010110010111100001000100101000011111011011001110110000100010111101",
   "11100101101001110000100111110011100101001101110011011100011100110101110001011100101",
   "11100101101001110000100111110011100101001101110011011100011100110101110001011100101",
   "11100101110000111110101001101100100010001010110111011010101101100100101010011100111",
   "11100101111000001100111000100111101110011110001100101011111010001001001000000110100",
   "11100101111000001100111000100111101110011110001100101011111010001001001000000110100",
   "11100101111111011011010100100101111001001101101110111101001111001101111110100100010",
   "11100110000110101001111101100111110001100011011001010000001010011010010101101001001",
   "11100110000110101001111101100111110001100011011001010000001010011010010101101001001",
   "11100110001101111000110011101110000110101101000110010111010000101101101111111010000",
   "11100110001101111000110011101110000110101101000110010111010000101101101111111010000",
   "11100110010101000111110110111001100111111100110001010011001001000001001100111100010",
   "11100110011100010111000111001011000100101000010101101111011010101101110010111011010",
   "11100110011100010111000111001011000100101000010101101111011010101101110010111011010",
   "11100110100011100110100100100011001100001001110000011111110000011001101011111101110",
   "11100110100011100110100100100011001100001001110000011111110000011001101011111101110",
   "11100110101010110110001111000010101101111110111111111100111110101100000011101101110",
   "11100110110010000110000110101010011001101010000100100010001111001000110001111111010",
   "11100110110010000110000110101010011001101010000100100010001111001000110001111111010",
   "11100110111001010110001011011010111110110001000001001010001111010100011111001000110",
   "11100110111001010110001011011010111110110001000001001010001111010100011111001000110",
   "11100111000000100110011101010101001100111101111011101100100100000001101111001011100",
   "11100111000111110110111100011001110011111110111101011011000000101000000000110000101",
   "11100111000111110110111100011001110011111110111101011011000000101000000000110000101",
   "11100111001111000111101000101001100011100110010011011111000010100101001101001011111",
   "11100111001111000111101000101001100011100110010011011111000010100101001101001011111",
   "11100111010110011000100010000101001011101010001111010111010001001010010110111001110",
   "11100111011101101001101000101101011100000101000111010101000001010100010011111011110",
   "11100111011101101001101000101101011100000101000111010101000001010100010011111011110",
   "11100111100100111010111100100011000100110101010110111001111101110001000001111011100",
   "11100111101100001100011101100110110101111101011111010101110011010010010001101001100",
   "11100111101100001100011101100110110101111101011111010101110011010010010001101001100",
   "11100111110011011110001011111001011111100100001000000100000001001110010111110001010",
   "11100111110011011110001011111001011111100100001000000100000001001110010111110001010",
   "11100111111010110000000111011011110001110011111111001001101110001111110001001011000",
   "11101000000010000010010000001110011100111011111001110011100001010100001000110111110",
   "11101000000010000010010000001110011100111011111001110011100001010100001000110111110",
   "11101000001001010100100110010010010001001110110100110011011110111011101101111111010",
   "11101000001001010100100110010010010001001110110100110011011110111011101101111111010",
   "11101000010000100111001001100111111111000011110100111111001010101001101000010010101",
   "11101000010111111001111010010000010110110110000111101101101100110101111001111011111",
   "11101000010111111001111010010000010110110110000111101101101100110101111001111011111",
   "11101000011111001100111000001100001001000101000011010101111100110001111101001111101",
   "11101000011111001100111000001100001001000101000011010101111100110001111101001111101",
   "11101000100110100000000011011100000110010100000111101100101111000000001101011100010",
   "11101000101101110011011100000000111111001010111110100011000111111111101001011111001",
   "11101000101101110011011100000000111111001010111110100011000111111111101001011111001",
   "11101000110101000111000001111011100100010101011100000100110011001100000000001100101",
   "11101000110101000111000001111011100100010101011100000100110011001100000000001100101",
   "11101000111100011010110101001100100110100011011111010110011110010011010101000111011",
   "11101001000011101110110101110100110110101001010010110100011001000001101101100110010",
   "11101001000011101110110101110100110110101001010010110100011001000001101101100110010",
   "11101001001011000011000011110101000101011111001100110000111001000011110101111000000",
   "11101001001011000011000011110101000101011111001100110000111001000011110101111000000",
   "11101001010010010111011111001110000100000001101111110011000010100001001101110111111",
   "11101001011001101100001000000000100011010001101011010101010100101110101101110100100",
   "11101001011001101100001000000000100011010001101011010101010100101110101101110100100",
   "11101001100001000000111110001101010100010011111100000100011011011010010010110000100",
   "11101001100001000000111110001101010100010011111100000100011011011010010010110000100",
   "11101001101000010110000001110101001000010001101100011110000100010000100011010000000",
   "11101001101111101011010010111000110000011000010101001111111000111100111100101111011",
   "11101001101111101011010010111000110000011000010101001111111000111100111100101111011",
   "11101001110111000000110001011000111101111001011101110110011101100101011010001000010",
   "11101001110111000000110001011000111101111001011101110110011101100101011010001000010",
   "11101001111110010110011101010110100010001010111100111100010011100010000100010110010",
   "11101001111110010110011101010110100010001010111100111100010011100010000100010110010",
   "11101010000101101100010110110010001110100110111000111001000000110001111101110010100",
   "11101010001101000010011101101100110100101011101000010000011011101101011001101100000",
   "11101010001101000010011101101100110100101011101000010000011011101101011001101100000",
   "11101010010100011000110010000111000101111011110010010001111011010110110000100111001",
   "11101010010100011000110010000111000101111011110010010001111011010110110000100111001",
   "11101010011011101111010100000001110011111110001111010111101100001010100011011101011",
   "11101010100011000110000011011101110000011110001001100110001001001111011110011110000",
   "11101010100011000110000011011101110000011110001001100110001001001111011110011110000",
   "11101010101010011101000000011011101101001010111101001011011010000111001101111001100",
   "11101010101010011101000000011011101101001010111101001011011010000111001101111001100",
   "11101010110001110100001010111100011011111000011000111110110101000000110110001101110",
   "11101010111001001011100011000000101110011110011111000000100101101101100001110001101",
   "11101010111001001011100011000000101110011110011111000000100101101101100001110001101",
   "11101011000000100011001000101001010110111001100100111001011000111000010110001000111",
   "11101011000000100011001000101001010110111001100100111001011000111000010110001000111",
   "11101011000111111010111011110111000111001010010100011010001100000010000011010011101",
   "11101011001111010010111100101010110001010101101011111100000010000001011111010110111",
   "11101011001111010010111100101010110001010101101011111100000010000001011111010110111",
   "11101011010110101011001011000101000111100100111110111111111100001001100001000100110",
   "11101011010110101011001011000101000111100100111110111111111100001001100001000100110",
   "11101011011110000011100111000110111100000101110110101110110111110101001100010111101",
   "11101011011110000011100111000110111100000101110110101110110111110101001100010111101",
   "11101011100101011100010000110001000001001010010010011001110000111011000011011010100",
   "11101011101100110101001000000100001001001000100111111001101000101000001111100101111",
   "11101011101100110101001000000100001001001000100111111001101000101000001111100101111",
   "11101011110100001110001101000001000110011011100100001111110001000100010101100000111",
   "11101011110100001110001101000001000110011011100100001111110001000100010101100000111",
   "11101011111011100111011111101000101011100010001100000101111101011110100111100010110",
   "11101100000011000000111111111011101010111111111100001110110111000101101010011001000",
   "11101100000011000000111111111011101010111111111100001110110111000101101010011001000",
   "11101100001010011010101101111010110111011100101010000110010110101001111111100001111",
   "11101100001010011010101101111010110111011100101010000110010110101001111111100001111",
   "11101100010001110100101001100111000011100100100100010010000010101100101001010110010",
   "11101100010001110100101001100111000011100100100100010010000010101100101001010110010",
   "11101100011001001110110011000001000010001000010011000001110010011010011101000111101",
   "11101100100000101001001010001001100101111100111000110000010101010100110111000000000",
   "11101100100000101001001010001001100101111100111000110000010101010100110111000000000",
   "11101100101000000011101111000001100001111011110010100011111111101001000100011111101",
   "11101100101000000011101111000001100001111011110010100011111111101001000100011111101",
   "11101100101111011110100001101001101001000010111000101111011011010110011001111100100",
   "11101100110110111001100010000010101110010100011111010010011110000100100111110001011",
   "11101100110110111001100010000010101110010100011111010010011110000100100111110001011",
   "11101100111110010100110000001101100100110111010110011011000011101011000100011000100",
   "11101100111110010100110000001101100100110111010110011011000011101011000100011000100",
   "11101101000101110000001100001010111111110110101011000110001101101001011111110100110",
   "11101101000101110000001100001010111111110110101011000110001101101001011111110100110",
   "11101101001101001011110101111011110010100010000111100001000111010011010110011010100",
   "11101101010100100111101101100000110000001101110011101010001110101110010111110000011",
   "11101101010100100111101101100000110000001101110011101010001110101110010111110000011",
   "11101101011100000011110010111010101100010010010101110010100010100101010111101110011",
   "11101101011100000011110010111010101100010010010101110010100010100101010111101110011",
   "11101101100011100000000110001010011010001100110010111110110100101111111111001100000",
   "11101101100011100000000110001010011010001100110010111110110100101111111111001100000",
   "11101101101010111100100111010000101101011110101111101001000001110000010010010110011",
   "11101101110010011001010110001110011001101110010000000001101101000111000010110101101",
   "11101101110010011001010110001110011001101110010000000001101101000111000010110101101",
   "11101101111001110110010011000100010010100101111000110001100010011111100011110011001",
   "11101101111001110110010011000100010010100101111000110001100010011111100011110011001",
   "11101110000001010011011101110011001011110100101111011010111011110011110110011011001",
   "11101110001000110000110110011011111001001110011010111011101100001010000101100001100",
   "11101110001000110000110110011011111001001110011010111011101100001010000101100001100",
   "11101110010000001110011100111111001110101011000100001110101111101100000110111100101",
   "11101110010000001110011100111111001110101011000100001110101111101100000110111100101",
   "11101110010111101100010001011110000000000111010110101110000000011001111001110011001",
   "11101110010111101100010001011110000000000111010110101110000000011001111001110011001",
   "11101110011111001010010011111001000001100100100000110100001111110111111000100100110",
   "11101110100110101000100100010001000111001000010100011111000101111001110110100011111",
   "11101110100110101000100100010001000111001000010100011111000101111001110110100011111",
   "11101110101110000111000010100111000100111101000111110001000100001011011111111101100",
   "11101110101110000111000010100111000100111101000111110001000100001011011111111101100",
   "11101110110101100101101110111011101111010001110101010011101110110111010100011010101",
   "11101110110101100101101110111011101111010001110101010011101110110111010100011010101",
   "11101110111101000100101001001111111010011001111100111001111010001100110011110001101",
   "11101111000100100011110001100100011010101101100100000001111101000110110101001000101",
   "11101111000100100011110001100100011010101101100100000001111101000110110101001000101",
   "11101111001100000011000111111010000100101001010110011000001000110011000000010101111",
   "11101111001100000011000111111010000100101001010110011000001000110011000000010101111",
   "11101111010011100010101100010001101100101110100110011001000101011011000010010110001",
   "11101111010011100010101100010001101100101110100110011001000101011011000010010110001",
   "11101111011011000010011110101100000111100011001101110100010011110000110100111110000",
   "11101111100010100010011111001010001001110001101110001110110011111110010010110101101",
   "11101111100010100010011111001010001001110001101110001110110011111110010010110101101",
   "11101111101010000010101101101100101000001001010001100101110001011001110000010111110",
   "11101111101010000010101101101100101000001001010001100101110001011001110000010111110",
   "11101111110001100011001010010100010111011101101010110001010011011111110010111111110",
   "11101111110001100011001010010100010111011101101010110001010011011111110010111111110",
   "11101111111001000011110101000010001100100111010110000111010011110011011111110100000",
   "11110000000000100100101101110110111100100011011001111110011001000101111011001110101",
   "11110000000000100100101101110110111100100011011001111110011001000101111011001110101",
   "11110000001000000101110100110011011100010011100111010000110111100101110011001110000",
   "11110000001000000101110100110011011100010011100111010000110111100101110011001110000",
   "11110000001111100111001001111000100000111110011001111111110110011000001110000010000",
   "11110000001111100111001001111000100000111110011001111111110110011000001110000010000",
   "11110000010111001000101101000110111111101110111001110110011001111011010111011001001",
   "11110000010111001000101101000110111111101110111001110110011001111011010111011001001",
   "11110000011110101010011110011111101101110100111010101100110011110100000110011011010",
   "11110000100110001100011110000011100000100100111101001011110111100111010110101100000",
   "11110000100110001100011110000011100000100100111101001011110111100111010110101100000",
   "11110000101101101110101011110011001101011000001111010000010101000000001110111001100",
   "11110000101101101110101011110011001101011000001111010000010101000000001110111001100",
   "11110000110101010001000111101111101001101100101100101110010111000011110000001100000",
   "11110000110101010001000111101111101001101100101100101110010111000011110000001100000",
   "11110000111100110011110001111001101011000100111111110101001000110011001000110001010",
   "11110001000100010110101010010010000111001000100001110010011110111101100101010010010",
   "11110001000100010110101010010010000111001000100001110010011110111101100101010010010",
   "11110001001011111001110000111001110011100011011011010110100111000010011100000100100",
   "11110001001011111001110000111001110011100011011011010110100111000010011100000100100",
   "11110001010011011101000101110001100110000110100101010111111011100100101101111110111",
   "11110001010011011101000101110001100110000110100101010111111011100100101101111110111",
   "11110001011011000000101000111010010100100111101001010110111101110000111000011101011",
   "11110001011011000000101000111010010100100111101001010110111101110000111000011101011",
   "11110001100010100100011010010100110101000001000010000010010100010101110100110001101",
   "11110001101010001000011010000001111101010001111011111010101111110010000000100101110",
   "11110001101010001000011010000001111101010001111011111010101111110010000000100101110",
   "11110001110001101100101000000010100011011110010101110111010011110101101100001000010",
   "11110001110001101100101000000010100011011110010101110111010011110101101100001000010",
   "11110001111001010001000100010111011101101111000001101001100110011011001010100000010",
   "11110001111001010001000100010111011101101111000001101001100110011011001010100000010",
   "11110010000000110101101111000001100010010001100100100010000011110110000000110110101",
   "11110010000000110101101111000001100010010001100100100010000011110110000000110110101",
   "11110010001000011010101000000001100111011000010111110100011000011010010001010000011",
   "11110010001111111111101111011000100011011010101001011011111111011100011110011110001",
   "11110010001111111111101111011000100011011010101001011011111111011100011110011110001",
   "11110010010111100101000101000111001100110100011100100000100111101011100101110101101",
   "11110010010111100101000101000111001100110100011100100000100111101011100101110101101",
   "11110010011111001010101001001110011010000110101001111010111101000101101100110100000",
   "11110010011111001010101001001110011010000110101001111010111101000101101100110100000",
   "11110010100110110000011011101111000001110111000000111001011000001000011111110110011",
   "11110010100110110000011011101111000001110111000000111001011000001000011111110110011",
   "11110010101110010110011100101001111010110000000111100100110010011110100000100001111",
   "11110010110101111100101011111111111011100001011011100101100001001010000001000000001",
   "11110010110101111100101011111111111011100001011011100101100001001010000001000000001",
   "11110010111101100011001001110001111010111111010010101000010100001110101011000110110",
   "11110010111101100011001001110001111010111111010010101000010100001110101011000110110",
   "11110011000101001001110110000000110000000010111011000011011011111010110001100101110",
   "11110011000101001001110110000000110000000010111011000011011011111010110001100101110",
   "11110011001100110000110000101101010001101010011100011011110011010001001010001101001",
   "11110011001100110000110000101101010001101010011100011011110011010001001010001101001",
   "11110011010100010111111001111000010110111000111000001010010000010100101111100011000",
   "11110011011011111111010001100010110110110110001010000000111001110110101001110001010",
   "11110011011011111111010001100010110110110110001010000000111001110110101001110001010",
   "11110011100011100110110111101101101000101111001000110000100010100111111101011110110",
   "11110011100011100110110111101101101000101111001000110000100010100111111101011110110",
   "11110011101011001110101100011001100011110101100110101110001010010000000000011000000",
   "11110011101011001110101100011001100011110101100110101110001010010000000000011000000",
   "11110011110010110110101111100111011111100000010010011000100011101000010011010010110",
   "11110011110010110110101111100111011111100000010010011000100011101000010011010010110",
   "11110011111010011111000001011000010011001010110110111110000000111111000001101011011",
   "11110100000010000111100001101100110110010101111101000010000101100001000110100101110",
   "11110100000010000111100001101100110110010101111101000010000101100001000110100101110",
   "11110100001001110000010000100110000000100111001011000011011100101100110111100101101",
   "11110100001001110000010000100110000000100111001011000011011100101100110111100101101",
   "11110100010001011001001110000100101001101001000110000001110111001110010110000110110",
   "11110100010001011001001110000100101001101001000110000001110111001110010110000110110",
   "11110100011001000010011010001001101001001011010010000100001101100110001000000011000",
   "11110100011001000010011010001001101001001011010010000100001101100110001000000011000",
   "11110100100000101011110100110101110111000010010010111110101000011011111000101001110",
   "11110100100000101011110100110101110111000010010010111110101000011011111000101001110",
   "11110100101000010101011110001010001011000111101100111000101110011101100010110001101",
   "11110100101111111111010110000111011101011010000100110011111000001100000110000001110",
   "11110100101111111111010110000111011101011010000100110011111000001100000110000001110",
   "11110100110111101001011100101110100101111101000001010001101001010111001000011010110",
   "11110100110111101001011100101110100101111101000001010001101001010111001000011010110",
   "11110100111111010011110010000000011100111001001010111010010000001000000110010100111",
   "11110100111111010011110010000000011100111001001010111010010000001000000110010100111",
   "11110101000110111110010101111101111010011100001101000011001001111110010010110110110",
   "11110101000110111110010101111101111010011100001101000011001001111110010010110110110",
   "11110101001110101001001000100111110110111000110110010101101110011100101010111000011",
   "11110101001110101001001000100111110110111000110110010101101110011100101010111000011",
   "11110101010110010100001001111111001010100110111001010101111111101010011101001111110",
   "11110101011101111111011010000100101110000011001101001001100000100111101010110111000",
   "11110101011101111111011010000100101110000011001101001001100000100111101010110111000",
   "11110101100101101010111000111001011001101111101101111110010001010110100001100101101",
   "11110101100101101010111000111001011001101111101101111110010001010110100001100101101",
   "11110101101101010110100110011110000110010011011101110001110000111010110101001000001",
   "11110101101101010110100110011110000110010011011101110001110000111010110101001000001",
   "11110101110101000010100010110011101100011010100100111000000101010000011001001100100",
   "11110101110101000010100010110011101100011010100100111000000101010000011001001100100",
   "11110101111100101110101101111011000100110110010010100011001000111001100000101011100",
   "11110101111100101110101101111011000100110110010010100011001000111001100000101011100",
   "11110110000100011011000111110101001000011100111101101001111110100110100101100000000",
   "11110110000100011011000111110101001000011100111101101001111110100110100101100000000",
   "11110110001100000111110000100010110000001010000101010000001010110111111101010010100",
   "11110110010011110100101000000100110100111110010001001101010011011010111111000101101",
   "11110110010011110100101000000100110100111110010001001101010011011010111111000101101",
   "11110110011011100001101110011100001111111111010010110100100100100011011110100111000",
   "11110110011011100001101110011100001111111111010010110100100100100011011110100111000",
   "11110110100011001111000011101001111010011000000101011100011100100010100001101110010",
   "11110110100011001111000011101001111010011000000101011100011100100010100001101110010",
   "11110110101010111100100111101110101101011000101111000110011100111011110101001000110",
   "11110110101010111100100111101110101101011000101111000110011100111011110101001000110",
   "11110110110010101010011010101011100010010110100001000111000001111010100101011100000",
   "11110110110010101010011010101011100010010110100001000111000001111010100101011100000",
   "11110110111010011000011100100001010010101011111000101101011111100111000001111000000",
   "11110110111010011000011100100001010010101011111000101101011111100111000001111000000",
   "11110111000010000110101101010000110111111000011111101100000101011101101110100001001",
   "11110111001001110101001100111011001011100001001101000000000111101001101011101000100",
   "11110111001001110101001100111011001011100001001101000000000111101001101011101000100",
   "11110111010001100011111011100001000111010000000101011010001110100010011000011000010",
   "11110111010001100011111011100001000111010000000101011010001110100010011000011000010",
   "11110111011001010010111001000011100100110100011100000110101100001110110111000111111",
   "11110111011001010010111001000011100100110100011100000110101100001110110111000111111",
   "11110111100001000010000101100011011110000010110011010101111000001110111001111011110",
   "11110111100001000010000101100011011110000010110011010101111000001110111001111011110",
   "11110111101000110001100001000001101100110100111101000100110001001011011110000001001",
   "11110111101000110001100001000001101100110100111101000100110001001011011110000001001",
   "11110111110000100001001011011111001011001001111011100101100100101111011101001001100",
   "11110111110000100001001011011111001011001001111011100101100100101111011101001001100",
   "11110111111000010001000100111100110011000110000010001000011101101001111100010010111",
   "11111000000000000001001101011011011110110010110101100100010111111010111110111110001",
   "11111000000000000001001101011011011110110010110101100100010111111010111110111110001",
   "11111000000111110001100100111100001000011111001100111111111011001100000111000001000",
   "11111000000111110001100100111100001000011111001100111111111011001100000111000001000",
   "11111000001111100010001011011111101010011111010010011010011011010101101000110000100",
   "11111000001111100010001011011111101010011111010010011010011011010101101000110000100",
   "11111000010111010011000001000110111111001100100011010100111111010001111011110010101",
   "11111000010111010011000001000110111111001100100011010100111111010001111011110010101",
   "11111000011111000100000101110011000001000101110001011011101101111111110000110000111",
   "11111000011111000100000101110011000001000101110001011011101101111111110000110000111",
   "11111000100110110101011001100100101010101111000011001111000001110100110100111001100",
   "11111000100110110101011001100100101010101111000011001111000001110100110100111001100",
   "11111000101110100110111100011100110110110001110100101101000010000001101100001000101",
   "11111000101110100110111100011100110110110001110100101101000010000001101100001000101",
   "11111000110110011000101110011100011111111100110111111011000010101000001011000101000",
   "11111000110110011000101110011100011111111100110111111011000010101000001011000101000",
   "11111000111110001010101111100100100001000100010101101111001010100101011010001001100",
   "11111001000101111100111111110101110101000001101110011010000000010000101011100110101",
   "11111001000101111100111111110101110101000001101110011010000000010000101011100110101",
   "11111001001101101111011111010001010110110011111010010000011100010000001110010010001",
   "11111001001101101111011111010001010110110011111010010000011100010000001110010010001",
   "11111001010101100010001101111000000001011111001010010101100010100101000111010010100",
   "11111001010101100010001101111000000001011111001010010101100010100101000111010010100",
   "11111001011101010101001011101010110000001101001001000100100010001111011100111011001",
   "11111001011101010101001011101010110000001101001001000100100010001111011100111011001",
   "11111001100101001000011000101010011110001100111010111010111011001011111101100011111",
   "11111001100101001000011000101010011110001100111010111010111011001011111101100011111",
   "11111001101100111011110100111000000110110010111111000010101010101100001101010100111",
   "11111001101100111011110100111000000110110010111111000010101010101100001101010100111",
   "11111001110100101111100000010100100101011001001111111100011110001010100101101110010",
   "11111001110100101111100000010100100101011001001111111100011110001010100101101110010",
   "11111001111100100011011011000000110101011111000100001010001100011011010010100110000",
   "11111001111100100011011011000000110101011111000100001010001100011011010010100110000",
   "11111010000100010111100100111101110010101001001110111001010101011011011000000010101",
   "11111010000100010111100100111101110010101001001110111001010101011011011000000010101",
   "11111010001100001011111110001100011000100010000000101101101000011111001101001110100",
   "11111010001100001011111110001100011000100010000000101101101000011111001101001110100",
   "11111010010100000000100110101101100010111001001000001011110001000001011000001010010",
   "11111010011011110101011110100010001101100011110010100100001001110011010110111010001",
   "11111010011011110101011110100010001101100011110010100100001001110011010110111010001",
   "11111010100011101010100101101011010100011100101100011101110110110001000010110110110",
   "11111010100011101010100101101011010100011100101100011101110110110001000010110110110",
   "11111010101011011111111100001001110011100100000010100001100101011000011010111100010",
   "11111010101011011111111100001001110011100100000010100001100101011000011010111100010",
   "11111010110011010101100001111110100110111111100010000100110011100110100010000010100",
   "11111010110011010101100001111110100110111111100010000100110011100110100010000010100",
   "11111010111011001011010111001010101010111010011001110100111101011010111110111001100",
   "11111010111011001011010111001010101010111010011001110100111101011010111110111001100",
   "11111011000011000001011011101110111011100101011010100010110001000011001011010110101",
   "11111011000011000001011011101110111011100101011010100010110001000011001011010110101",
   "11111011001010110111101111101100010101010110110111101101101001101110100000101110011",
   "11111011001010110111101111101100010101010110110111101101101001101110100000101110011",
   "11111011010010101110010011000011110100101010101000001111010001001100101111101001000",
   "11111011010010101110010011000011110100101010101000001111010001001100101111101001000",
   "11111011011010100101000101110110010110000010000111000111000111110111110001101111010",
   "11111011011010100101000101110110010110000010000111000111000111110111110001101111010",
   "11111011100010011100001000000100110110000100010100000110010011101010000011111111010",
   "11111011100010011100001000000100110110000100010100000110010011101010000011111111010",
   "11111011101010010011011001110000010001011101110100011011010101100010111000101000101",
   "11111011101010010011011001110000010001011101110100011011010101100010111000101000101",
   "11111011110010001010111010111001100101000000110011011110000101111001110000000001100",
   "11111011110010001010111010111001100101000000110011011110000101111001110000000001100",
   "11111011111010000010101011100001101101100101000011011011110111100010000111110101111",
   "11111100000001111010101011101001101000000111111110000011100001100000110000100100110",
   "11111100000001111010101011101001101000000111111110000011100001100000110000100100110",
   "11111100001001110010111011010010010001101100100101010001101111110011111001001111100",
   "11111100001001110010111011010010010001101100100101010001101111110011111001001111100",
   "11111100010001101011011010011100100111011011100011111101011010101111100001110001011",
   "11111100010001101011011010011100100111011011100011111101011010101111100001110001011",
   "11111100011001100100001001001001100110100011001110100100000101001111000100100100111",
   "11111100011001100100001001001001100110100011001110100100000101001111000100100100111",
   "11111100100001011101000111011010001100010111100011110110100001111101101000010000101",
   "11111100100001011101000111011010001100010111100011110110100001111101101000010000101",
   "11111100101001010110010101001111010110010010001101100101011111010110001010100100110",
   "11111100101001010110010101001111010110010010001101100101011111010110001010100100110",
   "11111100110001001111110010101010000001110010100001001110011010011100110110000100110",
   "11111100110001001111110010101010000001110010100001001110011010011100110110000100110",
   "11111100111001001001011111101011001100011101100000101000011000110010110100001010000",
   "11111100111001001001011111101011001100011101100000101000011000110010110100001010000",
   "11111101000001000011011100010011110011111101111010110001001001000101101101011101101",
   "11111101000001000011011100010011110011111101111010110001001001000101101101011101101",
   "11111101001000111101101000100100110110000100001100011010001010111100001010111010110",
   "11111101001000111101101000100100110110000100001100011010001010111100001010111010110",
   "11111101010000111000000100011111010000100110100000110101111101100000101001111010001",
   "11111101010000111000000100011111010000100110100000110101111101100000101001111010001",
   "11111101011000110010110000000100000001100000110010100101010101001011110110011011111",
   "11111101011000110010110000000100000001100000110010100101010101001011110110011011111",
   "11111101100000101101101011010100000110110100101100000100111000001111111110010100111",
   "11111101100000101101101011010100000110110100101100000100111000001111111110010100111",
   "11111101101000101000110110010000011110101001101000011010100010100110010000110111111",
   "11111101101000101000110110010000011110101001101000011010100010100110010000110111111",
   "11111101110000100100010000111010000111001100110100000011010000011111111110100100011",
   "11111101110000100100010000111010000111001100110100000011010000011111111110100100011",
   "11111101111000011111111011010001111110110001001101100000110000011100001100110111000",
   "11111101111000011111111011010001111110110001001101100000110000011100001100110111000",
   "11111110000000011011110101011001000011101111100110000111011100000011110010001001011",
   "11111110000000011011110101011001000011101111100110000111011100000011110010001001011",
   "11111110001000010111111111010000010100100110100010101100011000001100101110100100011",
   "11111110001000010111111111010000010100100110100010101100011000001100101110100100011",
   "11111110010000010100011000111000101111111010011100010011011100000110010110010100000",
   "11111110010000010100011000111000101111111010011100010011011100000110010110010100000",
   "11111110011000010001000010010011010100010101100000111101011111101111100010100101011",
   "11111110011000010001000010010011010100010101100000111101011111101111100010100101011",
   "11111110100000001101111011100001000000100111110100010110110001011000011110100101110",
   "11111110100000001101111011100001000000100111110100010110110001011000011110100101110",
   "11111110101000001011000100100010110011100111010000100101010010010001000110001100100",
   "11111110101000001011000100100010110011100111010000100101010010010001000110001100100",
   "11111110110000001000011101011001101100001111100110110111011010100101101100001101110",
   "11111110110000001000011101011001101100001111100110110111011010100101101100001101110",
   "11111110111000000110000110000110101001100010100000010010100100101010111110100101010",
   "11111110111000000110000110000110101001100010100000010010100100101010111110100101010",
   "11111111000000000011111110101010101010100111011110100001111111011010111110111100101",
   "11111111000000000011111110101010101010100111011110100001111111011010111110111100101",
   "11111111001000000010000111000110101110101011111100100101101000000100000110100001100",
   "11111111001000000010000111000110101110101011111100100101101000000100000110100001100",
   "11111111010000000000011111011011110101000011001111100001001011001011101100010100110",
   "11111111010000000000011111011011110101000011001111100001001011001011101100010100110",
   "11111111010111111111000111101010111101000110100111001011001101000101100101001110000",
   "11111111010111111111000111101010111101000110100111001011001101000101100101001110000",
   "11111111011111111101111111110101000110010101001110111100011001100001110101100001110",
   "11111111011111111101111111110101000110010101001110111100011001100001110101100001110",
   "11111111100111111101000111111011010000010100001110011110111010110010001100001100101",
   "11111111100111111101000111111011010000010100001110011110111010110010001100001100101",
   "11111111101111111100011111111110011010101110101010011101111000001000011111110110011",
   "11111111101111111100011111111110011010101110101010011101111000001000011111110110011",
   "11111111110111111100000111111111100101010101100101010100111011101111100110011000100",
      others => (others => '0'));
      	begin 
      return tmp;
      end init_rom;
	signal rom : memory_t := init_rom;
   signal Y0 :  std_logic_vector(82 downto 0);
begin
	process(clk)
   begin
   if(rising_edge(clk)) then
   	Y0 <= rom(  TO_INTEGER(unsigned(X))  );
   end if;
   end process;
    Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                              LogTable_1_9_74
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity LogTable_1_9_74 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(73 downto 0)   );
end entity;

architecture arch of LogTable_1_9_74 is
   -- Build a 2-D array type for the RoM
   subtype word_t is std_logic_vector(73 downto 0);
   type memory_t is array(0 to 511) of word_t;
   function init_rom
      return memory_t is 
      variable tmp : memory_t := (
   "00000000010000000000000000000011111111111111111110101010101010101011001011",
   "00000000110000000000000000000100000000000000000001010101010101010101110101",
   "00000001010000000000000000100100000000000000100100000000000000101000100000",
   "00000001110000000000000001100100000000000010100110101010101111100011001011",
   "00000010010000000000000011000100000000000111001001010101101000000101110110",
   "00000010110000000000000101000100000000001111001100000000110011010000100011",
   "00000011010000000000000111100100000000011011101110101100011101000011010011",
   "00000011110000000000001010100100000000101101110001011000110100011110000111",
   "00000100010000000000001110000100000001000110010100000110001011100001000101",
   "00000100110000000000010010000100000001100110010110110100110111001100010000",
   "00000101010000000000010110100100000010001110111001100101001111011111101110",
   "00000101110000000000011011100100000011000000111100010111101111011011100111",
   "00000110010000000000100001000100000011111101011111001100110101000000000101",
   "00000110110000000000100111000100000101000101100010000101000001001101010010",
   "00000111010000000000101101100100000110011010000101000000111000000011011101",
   "00000111110000000000110100100100000111111100001000000001000000100010110100",
   "00001000010000000000111100000100001001101100101011000110000100101011101011",
   "00001000110000000001000100000100001011101100101110010000110001011110010111",
   "00001001010000000001001100100100001101111101010001100001110110111011001111",
   "00001001110000000001010101100100010000011111010100111010001000000010101111",
   "00001010010000000001011111000100010011010011111000011010011010110101010110",
   "00001010110000000001101001000100010110011011111100000011101000010011100100",
   "00001011010000000001110011100100011001111000011111110110101100011110000000",
   "00001011110000000001111110100100011101101010100011110100100110010101010011",
   "00001100010000000010001010000100100001110011000111111110010111111010001010",
   "00001100110000000010010110000100100110010011001100010101000110001101010111",
   "00001101010000000010100010100100101011001011110000111001111001001111110000",
   "00001101110000000010101111100100110000011101110101101101111100000010010000",
   "00001110010000000010111101000100110110001010011010110010011100100101110110",
   "00001110110000000011001011000100111100010010100000001000101011111011100110",
   "00001111010000000011011001100101000010110111000101110001111110000100101010",
   "00001111110000000011101000100101001001111001001011101111101010000010010001",
   "00010000010000000011111000000101010001011001110010000011001001110101110000",
   "00010000110000000100001000000101011001011001111000101101111010100000011111",
   "00010001010000000100011000100101100001111010011111110001011100000100000000",
   "00010001110000000100101001100101101010111100100111001111010001100001111001",
   "00010010010000000100111011000101110100100001001111001001000000111011110110",
   "00010010110000000101001101000101111110101001010111100000010011010011101001",
   "00010011010000000101011111100110001001010110000000010110110100101011001101",
   "00010011110000000101110010100110010100101000001001101110010100000100100010",
   "00010100010000000110000110000110100000100000110011101000100011100001101111",
   "00010100110000000110011010000110101101000000111110000111011000000101000011",
   "00010101010000000110101110100110111010001001101001001100101001110000110100",
   "00010101110000000111000011100111000111111011110100111010010011100111100000",
   "00010110010000000111011001000111010110011000100001010010010011101011101011",
   "00010110110000000111101111000111100101100000101110010110101011000000000100",
   "00010111010000001000000101100111110101010101011100001001011101100111100001",
   "00010111110000001000011100101000000101110111101010101100110010100100111110",
   "00011000010000001000110100001000010111001000011010000010110011111011100010",
   "00011000110000001001001100001000101001001000101010001101101110101110011110",
   "00011001010000001001100100101000111011111001011011001111110011000001001000",
   "00011001110000001001111101101001001111011011101101001011010011110111000010",
   "00011010010000001010010111001001100011110000100000000010100111010011110110",
   "00011010110000001010110001001001111000111000110011111000000110011011011000",
   "00011011010000001011001011101010001110110101101000101110001101010001100111",
   "00011011110000001011100110101010100101100111111110100111011010111010101001",
   "00011100010000001100000010001010111101010000110101100110010001011010110000",
   "00011100110000001100011110001011010101110001001101101101010101110110010111",
   "00011101010000001100111010101011101111001010000110111111010000010010000101",
   "00011101110000001101010111101100001001011100100001011110101011110010101010",
   "00011110010000001101110101001100100100101001011101001110010110011101000011",
   "00011110110000001110010011001101000000110001111010010001000001010110010101",
   "00011111010000001110110001101101011101110110111000101001100000100011110010",
   "00011111110000001111010000101101111011111001011000011010101011001010110111",
   "00100000010000001111110000001110011010111010011001100111011011010001001100",
   "00100000110000010000010000001110111010111010111100010010101101111100100111",
   "00100001010000010000110000101111011011111100000000011111100011010011000111",
   "00100001110000010001010001101111111101111110100110010000111110011010111000",
   "00100010010000010001110011010000100001000011101101101010000101011010010011",
   "00100010110000010010010101010001000101001100010110101110000001010111111110",
   "00100011010000010010110111110001101010011001100001011111111110011010101000",
   "00100011110000010011011010110010010000101100001110000011001011101001010010",
   "00100100010000010011111110010010111000000101011100011010111011001011000111",
   "00100100110000010100100010010011100000100110001100101010100010000111100000",
   "00100101010000010101000110110100001010001111011110110101011000100110000010",
   "00100101110000010101101011110100110101000010010010111110111001101110100011",
   "00100110010000010110010001010101100000111111101001001010100011101001000010",
   "00100110110000010110110111010110001110001000100001011011110111011101110001",
   "00100111010000010111011101110110111100011101111011110110011001010101001101",
   "00100111110000011000000100110111101100000000111000011101110000011000000010",
   "00101000010000011000101100011000011100110010010111010101100110101111001010",
   "00101000110000011001010100011001001110110011011000100001101001100011101111",
   "00101001010000011001111100111010000010000100111100000101101000111111001010",
   "00101001110000011010100101111010110110101000000010000101011000001011000010",
   "00101010010000011011001111011011101100011101101010100100101101010001001101",
   "00101010110000011011111001011100100011100110110101100111100001011011110010",
   "00101011010000011100100011111101011100000100100011010001110000110101000110",
   "00101011110000011101001110111110010101110111110011100111011010100111110000",
   "00101100010000011101111010011111010001000001100110101100100000111110100101",
   "00101100110000011110100110100000001101100010111100100101001001000100101100",
   "00101101010000011111010011000001001011011100110101010101011011000101011010",
   "00101101110000100000000000000010001010110000010001000001100010001100010110",
   "00101110010000100000101101100011001011011110001111101101101100100101011001",
   "00101110110000100001011011100100001101100111110001011110001011011100101011",
   "00101111010000100010001010000101010001001101110110010111010010111110100110",
   "00101111110000100010111001000110010110010001011110011101011010010111110111",
   "00110000010000100011101000100111011100110011101001110100111011110101011000",
   "00110000110000100100011000101000100100110101011000100010010100100100011010",
   "00110001010000100101001001001001101110010111101010101010000100110010011100",
   "00110001110000100101111010001010111001011011100000010000101111101101010010",
   "00110010010000100110101011101100000110000001111001011010111011100011000000",
   "00110010110000100111011101101101010100001011110110001101010001100001111110",
   "00110011010000101000010000001110100011111010010110101100011101111000110110",
   "00110011110000101001000011001111110101001110011010111101001111110110100101",
   "00110100010000101001110110110001001000001001000011000100011001101010011010",
   "00110100110000101010101010110010011100101011001111000110110000100011111010",
   "00110101010000101011011111010011110010110101111111001001001100110010111010",
   "00110101110000101100010100010101001010101010010011010000101001100111100110",
   "00110110010000101101001001110110100100001001001011100010000101010010011011",
   "00110110110000101101111111110111111111010011101000000010100001000100001100",
   "00110111010000101110110110011001011100001010101000110111000001001101111110",
   "00110111110000101111101101011010111010101111001110000100101101000001001100",
   "00111000010000110000100100111100011011000010010111110000101110101111100110",
   "00111000110000110001011100111101111101000101000110000000010011101011001111",
   "00111001010000110010010101011111100000111000011000111000101100000110100000",
   "00111001110000110011001110100001000110011101010000011111001011010100001000",
   "00111010010000110100001000000010101101110100101100111001000111100111001001",
   "00111010110000110101000010000100010110111111101110001011111010010010111100",
   "00111011010000110101111100100110000001111111010100011100111111101011010001",
   "00111011110000110110110111100111101110110100011111110001110111000100001010",
   "00111100010000110111110011001001011101100000010000010000000010110010000011",
   "00111100110000111000101111001011001110000011100101111101001000001001101100",
   "00111101010000111001101011101101000000011111100000111110101111100000001100",
   "00111101110000111010101000101110110100110101000001011010100100001011000000",
   "00111110010000111011100110010000101011000101000111010110010100011111111111",
   "00111110110000111100100100010010100011010000110010110111110001110101010010",
   "00111111010000111101100010110100011101011001000100000100110000100001011100",
   "00111111110000111110100001110110011001011110111011000011000111111011011000",
   "01000000010000111111100001011000010111100011010111111000110010011010010110",
   "01000000110001000000100001011010010111100111011010101011101101010110000010",
   "01000001010001000001100001111100011001101100000011100001111001000110011010",
   "01000001110001000010100010111110011101110010010010100001011001000011111010",
   "01000010010001000011100100100000100011111011000111110000010011100111010011",
   "01000010110001000100100110100010101100000111100011010100110010001001101111",
   "01000011010001000101101001000100110110011000100101010101000001000100110000",
   "01000011110001000110101100000111000010101111001101110111001111110010010100",
   "01000100010001000111101111101001010001001100011101000001110000101100101110",
   "01000100110001001000110011101011100001110001010010111010111001001110101100",
   "01000101010001001001111000001101110100011110101111101001000001110011010110",
   "01000101110001001010111101010000001001010101110011010010100101110110001110",
   "01000110010001001100000010110010100000010111011101111110000011110011001110",
   "01000110110001001101001000110100111001100100101111110001111101000110101010",
   "01000111010001001110001111010111010100111110101000110100110110001101010100",
   "01000111110001001111010110011001110010100110001001001101010110100100010011",
   "01001000010001010000011101111100010010011100010001000010001000101001001100",
   "01001000110001010001100101111110110100100010000000011001111001111001111110",
   "01001001010001010010101110100001011000111000010111011011011010110101000011",
   "01001001110001010011110111100011111111100000010110001101011110111001010000",
   "01001010010001010101000001000110101000011010111100110110111100100101110100",
   "01001010110001010110001011001001010011101001001011011110101101011010011011",
   "01001011010001010111010101101100000001001100000010001011101101110111001110",
   "01001011110001011000100000101110110001000100100001000100111101011100101111",
   "01001100010001011001101100010001100011010011101000010001011110101011111110",
   "01001100110001011010111000010100010111111010010111111000010111000110010110",
   "01001101010001011100000100110111001110111001110000000000101111001101110000",
   "01001101110001011101010001111010001000010010110000110001110010100100100001",
   "01001110010001011110011111011101000100000110011010010010101111101101011010",
   "01001110110001011111101101100000000010010101101100101010111000001011101000",
   "01001111010001100000111100000011000011000001101000000001100000100010111010",
   "01001111110001100010001011000110000110001011001100011110000000010111010110",
   "01010000010001100011011010101001001011110011011010000111110010001101100101",
   "01010000110001100100101010101100010011111011010001000110010011101010101011",
   "01010001010001100101111011001111011110100011110001100001000101010100001010",
   "01010001110001100111001100010010101011101101111011011111101010110000000010",
   "01010010010001101000011101110101111011011010101111001001101010100100110100",
   "01010010110001101001101111111001001101101011001100100110101110011001011100",
   "01010011010001101011000010011100100010100000010011111110100010110101010110",
   "01010011110001101100010101011111111001111011000101011000110111100000011101",
   "01010100010001101101101001000011010011111100100000111101011111000011001100",
   "01010100110001101110111101000110110000100101100110110100001111000110011100",
   "01010101010001110000010001101010001111110111010111000101000000010011100110",
   "01010101110001110001100110101101110001110010110001110111101110010100100010",
   "01010110010001110010111100010001010110011000110111010100010111110011101000",
   "01010110110001110100010010010100111101101010100111100010111110011011110010",
   "01010111010001110101101000111000100111101001000010101011100110111000011000",
   "01010111110001110110111111111100010100010101001000110110011000110101010001",
   "01011000010001111000010111100000000011101111111010001011011110111110111001",
   "01011000110001111001101111100011110101111010010110110011000111000010001001",
   "01011001010001111011001000000111101010110101011110110101100001101100011100",
   "01011001110001111100100001001011100010100010010010011011000010101011110000",
   "01011010010001111101111010101111011101000001110001101100000000101110100010",
   "01011010110001111111010100110011011010010100111100110000110101100011110000",
   "01011011010010000000101111010111011010011100110011110001111101111010111101",
   "01011011110010000010001010011011011101011010010110110111111001100100001010",
   "01011100010010000011100101111111100011001110100110001011001011001111111110",
   "01011100110010000101000010000011101011111010100001110100011000101111100000",
   "01011101010010000110011110100111110111011111001001111100001010110100011000",
   "01011101110010000111111011101100000101111101011110101011001101010000110010",
   "01011110010010001001011001010000010111010110100000001010001110110111100001",
   "01011110110010001010110111010100101011101011001110100010000001011011110100",
   "01011111010010001100010101111001000010111100101001111011011001110001100001",
   "01011111110010001101110100111101011101001011110010011111001111101101000010",
   "01100000010010001111010100100001111010011001101000010110011110000011010010",
   "01100000110010010000110100100110011010100111001011101010000010101001110011",
   "01100001010010010010010101001010111101110101011100100010111110010110101000",
   "01100001110010010011110110001111100100000101011011001010010101000000011010",
   "01100010010010010101010111110100001101011000000111101001001101011110010100",
   "01100010110010010110111001111000111001101110100010001000110001101000001010",
   "01100011010010011000011100011101101001001001101010110010001110010110010000",
   "01100011110010011001111111100010011011101010100001101110110011100001100011",
   "01100100010010011011100011000111010001010010000111000111110100000011100001",
   "01100100110010011101000111001100001010000001011011000110100101110110010000",
   "01100101010010011110101011110001000101111001011101110100100001110100011100",
   "01100101110010100000010000110110000100111011001111011011000011111001010010",
   "01100110010010100001110110011011000111000111110000000011101011000000101100",
   "01100110110010100011011100100000001100011111111111110111111001000111000110",
   "01100111010010100101000011000101010101000100111111000001010011001001100000",
   "01100111110010100110101010001010100000110111101101101001100001000101100110",
   "01101000010010101000010001101111101111111001001011111010001101111001100100",
   "01101000110010101001111001110101000010001010011001111101000111100100010100",
   "01101001010010101011100010011010010111101100010111111011111111000101010010",
   "01101001110010101101001011011111110000100000000110000000101000011100100100",
   "01101010010010101110110101000101001100100110100100010100111010101010110010",
   "01101010110010110000011111001010101100000000110011000010101111110001010100",
   "01101011010010110010001001110000001110101111110010010100000100110010000010",
   "01101011110010110011110100110101110100110100100010010010111001101111100000",
   "01101100010010110101100000011011011110010000000011001001010001101100111010",
   "01101100110010110111001100100001001011000011010101000001010010101110000100",
   "01101101010010111000111001000110111011001111011000000101000101110111011000",
   "01101101110010111010100110001100101110110101001100011110110111001101111101",
   "01101110010010111100010011110010100101110101110010011000110101110111011110",
   "01101110110010111110000001111000100000010010001001111101010011111010010100",
   "01101111010010111111110000011110011110001011010011010110100110011101011110",
   "01101111110011000001011111100100011111100010001110101111000101101000100110",
   "01110000010011000011001111001010100100010111111100010001001100100011111101",
   "01110000110011000100111111010000101100101101011100000111011001011000100010",
   "01110001010011000110101111110110111000100011101110011100001101001111111010",
   "01110001110011001000100000111101000111111011110011011010001100010100010110",
   "01110010010011001010010010100011011010110110101011001011111101110000110010",
   "01110010110011001100000100101001110001010101010101111100001011110000110100",
   "01110011010011001101110111010000001011011000110011110101100011100000101101",
   "01110011110011001111101010010110101001000010000101000010110101001101011000",
   "01110100010011010001011101111101001010010010001001101110110100000100011010",
   "01110100110011010011010010000011101111001010000010000100010110010100001000",
   "01110101010011010101000110101010010111101010101110001110010101001011011101",
   "01110101110011010110111011110001000011110101001110010111101100111010000100",
   "01110110010011011000110001010111110011101010100010101011011100110000010000",
   "01110110110011011010100111011110100111001011101011010100100110111111000100",
   "01110111010011011100011110000101011110011001101000011110010000111000001101",
   "01110111110011011110010101001100011001010101011010010011100010101110000100",
   "01111000010011100000001100110011011000000000000000111111100111110011110000",
   "01111000110011100010000100111010011010011010011100101101101110011101000100",
   "01111001010011100011111101100001100000100101101101101001000111111110100001",
   "01111001110011100101110110101000101010100010110011111101001000101101010100",
   "01111010010011100111110000001111111000010010101111110101000111111111010111",
   "01111010110011101001101010010111001001110110100001011100100000001011010100",
   "01111011010011101011100100111110011111001111001000111110101110101000100000",
   "01111011110011101101100000000101111000011101100110100111010011101111000000",
   "01111100010011101111011011101101010101100010111010100001110010110111100101",
   "01111100110011110001010111110100110110100000000100111001110010011011110001",
   "01111101010011110011010100011100011011010110000101111010111011110101110010",
   "01111101110011110101010001100100000100000101111101110000111011100000100111",
   "01111110010011110111001111001011110000110000101100100111100000110111111100",
   "01111110110011111001001101010011100001010111010010101010011110011000001110",
   "01111111010011111011001011111011010101111010110000000101101001011110100110",
   "01111111110011111101001011000011001110011100000101000100111010101000111111",
   "10000000000011111110001010110011001100001100010000011101110011111101110000",
   "10000000100100000000001010101011001010101100010001001001100110101011111010",
   "10000001000100000010001011000011001101001100101001110111011001110100001000",
   "10000001100100000100001011111011010011101110011010110011010000010110111110",
   "10000010000100000110001101010011011110010010100100001001010000010101101101",
   "10000010100100001000001111001011101100111010000110000101100010110010011000",
   "10000011000100001010010001100011111111100110000000110100010011101111110011",
   "10000011100100001100010100011100010110010111010100100001110010010001100010",
   "10000100000100001110010111110100110001001111000001011010010000011011111100",
   "10000100100100010000011011101101010000001110000111101010000011010100000101",
   "10000101000100010010100000000101110011010101100111011101100010111111111000",
   "10000101100100010100100100111110011010100110100001000001001010100101111101",
   "10000110000100010110101010010111000110000001110100100001011000001101110001",
   "10000110100100011000110000001111110101101000100010001010101100111111100001",
   "10000111000100011010110110101000101001011011101010001001101101000100001100",
   "10000111100100011100111101100001100001011100001100101010111111100101100110",
   "10001000000100011111000100111010011101101011001001111011001110101110010010",
   "10001000100100100001001100110011011110001001100010000111000111101001101001",
   "10001001000100100011010101001100100010111000010101011011011010100011110101",
   "10001001100100100101011110000101101011111000100100000100111010101001110011",
   "10001010000100100111100111011110111001001011001110010000011110001001010101",
   "10001010100100101001110001011000001010110001010100001010111110010000111110",
   "10001011000100101011111011110001100000101011110110000001010111010000001000",
   "10001011100100101110000110101010111010111011110100000000101000010110111110",
   "10001100000100110000010010000100011001100010001110010101110011110110100000",
   "10001100100100110010011101111101111100100000000101001101111111000000100011",
   "10001101000100110100101010010111100011110110011000110110010010000111101111",
   "10001101100100110110110111010001001111100110001001011011111000011111100011",
   "10001110000100111001000100101010111111110000010111001100000000011100001111",
   "10001110100100111011010010100100110100010110000010010011111011010010111100",
   "10001111000100111101100000111110101101011000001011000000111101011001100110",
   "10001111100100111111101111111000101010110111110001100000011110000111000000",
   "10010000000101000001111111010010101100110101110101111111110111110010101111",
   "10010000100101000100001111001100110011010011011000101100100111110101010011",
   "10010001000101000110011111100110111110010001011001110100001110100111111101",
   "10010001100101001000110000100001001101110000111001100100001111100100111000",
   "10010010000101001011000001111011100001110010111000001010010001000111000011",
   "10010010100101001101010011110101111010011000010101110011111100101010010101",
   "10010011000101001111100110010000010111100010010010101110111110101011011001",
   "10010011100101010001111001001010111001010001101111001001000110100111110101",
   "10010100000101010100001100100101011111100111101011010000000110111110000011",
   "10010100100101010110100000100000001010100101000111010001110101001101010110",
   "10010101000101011000110100111010111010001011000011011100001001110101110110",
   "10010101100101011011001001110101101110011010011111111101000000011000100110",
   "10010110000101011101011111010000100111010100011101000010010111010111011111",
   "10010110100101011111110101001011100100111001111010111010010000010101010010",
   "10010111000101100010001011100110100111001011111001110010101111110101101000",
   "10010111100101100100100010100001101110001011011001111001111101011101000011",
   "10011000000101100110111001111100111001111001011011011110000011110000111101",
   "10011000100101101001010001111000001010010110111110101101010000010111101011",
   "10011001000101101011101010010011011111100101000011110101110011111000011000",
   "10011001100101101110000011001110111001100100101011000110000001111011001010",
   "10011010000101110000011100101010011000010110110100101100010001001000111111",
   "10011010100101110010110110100101111011111100100000110110111011001011101111",
   "10011011000101110101010001000001100100010110101111110100011100101110001110",
   "10011011100101110111101011111101010001100110100001110011010101011100000110",
   "10011100000101111010000111011001000011101100110111000010001000000001111110",
   "10011100100101111100100011010100111010101010101111101111011010001101010101",
   "10011101000101111110111111110000110110100001001100001001110100101100101000",
   "10011101100110000001011100101100110111010001001100100000000011001111001011",
   "10011110000110000011111010001000111100111011110001000000110100100101001111",
   "10011110100110000110011000000101000111100001111001111010111010011111111111",
   "10011111000110001000110110100001010111000100100111011101001001110001100011",
   "10011111100110001011010101011101101011100100111001110110011010001100111011",
   "10100000000110001101110100111010000101000011110001010101100110100110000110",
   "10100000100110010000010100110110100011100010001110001001101100110001111101",
   "10100001000110010010110101010011000111000001010000100001101101100110010110",
   "10100001100110010101010110001111101111100001111000101100101100111010000011",
   "10100010000110010111110111101100011101000101000110111001110001100100110001",
   "10100010100110011010011001101001001111101011111011011000000101011111001011",
   "10100011000110011100111100000110000111010111010110010110110101100010111001",
   "10100011100110011111011111000011000100001000011000000101010001101010011111",
   "10100100000110100010000010100000000110000000000000110010101100110001011110",
   "10100100100110100100100110011101001100111111010000101110011100110100010110",
   "10100101000110100111001010111010011001000111001000000111111010110000100010",
   "10100101100110101001101111110111101010011000100111001110100010100100011100",
   "10100110000110101100010101010101000000110100101110010001110011001111011101",
   "10100110100110101110111011010010011100011100011101100001001110110001111010",
   "10100111000110110001100001101111111101010000110101001100011010001101000111",
   "10100111100110110100001000101101100011010010110101100010111101100011010111",
   "10101000000110110110110000001011001110100011011110110100100011110111111011",
   "10101000100110111001011000001000111111000011110001010000111011001111000100",
   "10101001000110111100000000100110110100110100101101000111110100101110000000",
   "10101001100110111110101001100100101111110111010010101001000100011010111110",
   "10101010000111000001010011000010110000001100100010000100100001011101001011",
   "10101010100111000011111101000000110101110101011011101010000101111100110101",
   "10101011000111000110100111011111000000110010111111101001101111000011001001",
   "10101011100111001001010010011101010001000110001110010011011100111010010011",
   "10101100000111001011111101111011100110110000000111110111010010101101100010",
   "10101100100111001110101001111010000001110001101100100101010110101001000001",
   "10101101000111010001010110011000100010001011111100101101110001111010000000",
   "10101101100111010100000011010111000111111111111000100000110000101110101101",
   "10101110000111010110110000110101110011001110100000001110100010010110011000",
   "10101110100111011001011110110100100011111000110100000111011001000001010001",
   "10101111000111011100001101010011011001111111110100011011101010000000101010",
   "10101111100111011110111100010010010101100100100001011011101101100110111000",
   "10110000000111100001101011110001010110100111111011010111111111000111001110",
   "10110000100111100100011011110000011101001011000010100000111100110110000100",
   "10110001000111100111001100001111101001001110110111000111001000001000110011",
   "10110001100111101001111101001110111010110100011001011011000101010101110110",
   "10110010000111101100101110101110010001111100101001101101011011110100101011",
   "10110010100111101111100000101101101110101000101000001110110101111101110010",
   "10110011000111110010010011001101010000111001010101010000000001001010101101",
   "10110011100111110101000110001100111000101111110001000001101101110110000100",
   "10110100000111110111111001101100100110001100111011110100101111011011011110",
   "10110100100111111010101101101100011001010001110101111001111100010111101001",
   "10110101000111111101100010001100010001111111011111100010001110001000010101",
   "10110101101000000000010111001100010000010110111000111110100001001100010101",
   "10110110001000000011001100101100010100011001000010011111110101000011100001",
   "10110110101000000110000010101100011110000110111100010111001100001110110101",
   "10110111001000001000111001001100101101100001100110110101101100010000010001",
   "10110111101000001011110000001101000010101010000010001100011101101010111010",
   "10111000001000001110100111101101011101100001001110101100101100000010111000",
   "10111000101000010001011111101101111110001000001100100111100101111101011011",
   "10111001001000010100011000001110100100011111111100001110011101000000110100",
   "10111001101000010111010001001111010000101001011101110010100101110100011110",
   "10111010001000011010001010110000000010100101110001100101011000000000110101",
   "10111010101000011101000100110000111010010101110111111000001110001111011100",
   "10111011001000011111111111010001110111111010110000111100100110001010111111",
   "10111011101000100010111010010010111011010101011101000100000000011111001010",
   "10111100001000100101110101110100000100100110111100100000000000111000110101",
   "10111100101000101000110001110101010011110000001111100010001110000101111011",
   "10111101001000101011101110010110101000110010010110011100010001110101011110",
   "10111101101000101110101011011000000011101110010001011111111000110111101000",
   "10111110001000110001101000111001100100100101000000111110110010111101101000",
   "10111110101000110100100110111011001011010111100101001010110010111001110110",
   "10111111001000110111100101011100111000000110111110010101101110011111110001",
   "10111111101000111010100100011110101010110100001100110001011110100011111110",
   "11000000001000111101100100000000100011100000010000101111111110111100001011",
   "11000000101001000000100100000010100010001100001010100011001110011111001111",
   "11000001001001000011100100100100100110111000111010011101001111000101000110",
   "11000001101001000110100101100110110001100111100000110000000101100110110111",
   "11000010001001001001100111001001000010011000111101101101111001111110110000",
   "11000010101001001100101001001011011001001110010001101000110111001000001000",
   "11000011001001001111101011101101110110001000011100110011001010111111100000",
   "11000011101001010010101110110000011001001000011111011111000110100010100000",
   "11000100001001010101110010010011000010001111011001111110111101101111111010",
   "11000100101001011000110110010101110001011110001100100101000111100111101010",
   "11000101001001011011111010111000100110110101110111100011111110001010110101",
   "11000101101001011110111111111011100010010111011011001101111110011011101010",
   "11000110001001100010000101011110100100000011110111110101101000011101100010",
   "11000110101001100101001011100001101011111100001101101101011111010100111111",
   "11000111001001101000010010000100111010000001011101001000001001000111110000",
   "11000111101001101011011001001000001110010100100110011000001110111100101100",
   "11001000001001101110100000101011101000110110101001110000011100111011110110",
   "11001000101001110001101000101111001001101000100111100011100010001110011100",
   "11001001001001110100110001010010110000101011100000000100010000111110110101",
   "11001001101001110111111010010110011110000000010011100101011110011000100110",
   "11001010001001111011000011111010010001101000000010011010000010101000011110",
   "11001010101001111110001101111110001011100011101100110100111000111100011001",
   "11001011001010000001011000100010001011110100010011001000111111100011011101",
   "11001011101010000100100011100110010010011010110101101001010111101101111101",
   "11001100001010000111101111001010011111011000010100101001000101101101011001",
   "11001100101010001010111011001110110010101101110000011011010000110100011100",
   "11001101001010001110000111110011001100011100001001010011000011010110111110",
   "11001101101010010001010100110111101100100100011111100011101010101010000100",
   "11001110001010010100100010011100010011000111110011100000010111000100000001",
   "11001110101010010111110000100001000000000111000101011100011011111100010011",
   "11001111001010011010111111000101110011100011010101101011001111101011100111",
   "11001111101010011110001110001010101101011101100100100000001011101011110111",
   "11010000001010100001011101101111101101110110110010001110101100011000001100",
   "11010000101010100100101101110100110100101111111111001010010001001100111010",
   "11010001001010100111111110011010000010001010001011100110011100100111100110",
   "11010001101010101011001111011111010110000110010111110110110100000111000001",
   "11010010001010101110100001000100110000100101100100001111000000001011001110",
   "11010010101010110001110011001010010001101000110001000010101100010101011010",
   "11010011001010110101000101101111111001010000111110100101100111001000000101",
   "11010011101010111000011000110101100111011111001101001011100010000110111011",
   "11010100001010111011101100011011011100010100011101001000010001110110111010",
   "11010100101010111111000000100001010111110001101110101111101101111110001101",
   "11010101001011000010010101000111011001111000000010010101110001000100010000",
   "11010101101011000101101010001101100010101000011000001110011000110001101110",
   "11010110001011001000111111110011110010000011110000101101100101110000100011",
   "11010110101011001100010101111010001000001011001100000111011011101011111011",
   "11010111001011001111101100100000100100111111101010110000000001010000010010",
   "11010111101011010011000011100111001000100010001100111011100000001011010101",
   "11011000001011010110011011001101110010110011110010111110000101001100000000",
   "11011000101011011001110011010100100011110101011101001100000000000010100011",
   "11011001001011011101001011111011011011101000001011111001100011100000011101",
   "11011001101011100000100101000010011010001100111111011011000101011000011110",
   "11011010001011100011111110101001011111100100111000000100111110011110101010",
   "11011010101011100111011000110000101011110000110110001011101010101000010100",
   "11011011001011101010110011010111111110110001111010000011101000101100000010",
   "11011011101011101110001110011111011000101001000100000001011010100001101101",
   "11011100001011110001101010000110111001010111010100011001100101000010011111",
   "11011100101011110101000110001110100000111101101011100000110000001000110100",
   "11011101001011111000100010110110001111011101001001101011100110110000011101",
   "11011101101011111011111111111110000100110110101111001110110110110110011011",
   "11011110001011111111011101100110000001001011011100011111010001011001000101",
   "11011110101100000010111011101110000100011100010001110001101010011000000010",
   "11011111001100000110011010010110001110101010001111011010111000110100001111",
   "11011111101100001001111001011110011111110110010101101111110110101111111011",
   "11100000001100001101011001000110111000000001100101000101100001001110101010",
   "11100000101100010000111001001111010111001100111101110000111000010101010100",
   "11100001001100010100011001110111111101011001100000000110111111001010000011",
   "11100001101100010111111011000000101010101000001100011100111011110100011000",
   "11100010001100011011011100101001011110111010000011000111110111011101001000",
   "11100010101100011110111110110010011010010000000100011100111110001110011011",
   "11100011001100100010100001011011011100101011010000110001011111010011101111",
   "11100011101100100110000100100100100110001100101000011010101100111001111001",
   "11100100001100101001101000001101110110110101001011101101111100001111000001",
   "11100100101100101101001100010111001110100101111011000000100101100010100100",
   "11100101001100110000110001000000101101011111110110101000000100000101010110",
   "11100101101100110100010110001010010011100011111110111001110110001001100010",
   "11100110001100110111111011110100000000110011010100001011011101000010100111",
   "11100110101100111011100001111101110101001110110110110010011101000101011010",
   "11100111001100111111001000100111110000110111100111000100011101101000001001",
   "11100111101101000010101111110001110011101110100101010111001001000010010110",
   "11101000001101000110010111011011111101110100110010000000001100101100111011",
   "11101000101101001001111111100110001111001011001101010101011001000010001001",
   "11101001001101001101101000010000100111110010110111101100100001011101101000",
   "11101001101101010001010001011011000111101100110001011011011100011100011000",
   "11101010001101010100111011000101101110111001111010111000000011011100101111",
   "11101010101101011000100101010000011101011011010100011000010010111110011100",
   "11101011001101011100001111111011010011010001111110010010001010100010100110",
   "11101011101101011111111011000110010000011110111000111011101100101011101101",
   "11101100001101100011100110110001010101000011000100101010111110111101100110",
   "11101100101101100111010010111100100000111111100001110110001001111101100010",
   "11101101001101101010111111100111110100010101010000110011011001010010001001",
   "11101101101101101110101100110011001111000101010001111000111011100011011101",
   "11101110001101110010011010011110110001010000100101011101000010011010111000",
   "11101110101101110110001000101010011010111000001011110110000010100011001110",
   "11101111001101111001110111010110001011111101000101011010010011101000101100",
   "11101111101101111101100110100010000100100000010010100000010000011000111001",
   "11110000001110000001010110001110000100100010110011011110010110100010110101",
   "11110000101110000101000110011010001100000101101000101011000110110110111011",
   "11110001001110001000110111000110011011001001110010011101000101000111000000",
   "11110001101110001100101000010010110001110000010001001010111000000110010100",
   "11110010001110010000011001111111001111111010000101001011001001101001100000",
   "11110010101110010100001100001011110101101000001110110100100110100110101001",
   "11110011001110010111111110111000100010111011101110011101111110110101001111",
   "11110011101110011011110010000101010111110101100100011110000101001110001101",
   "11110100001110011111100101110010010100010110110001001011101111101011111001",
   "11110100101110100011011001111111011000100000010100111101110111001010000101",
   "11110101001110100111001110101100100100010011010000001011010111100101111110",
   "11110101101110101011000011111001110111110000100011001011001111111110001111",
   "11110110001110101110111001100111010010111001001110010100100010010010111011",
   "11110110101110110010101111110100110101101110010001111110010011100101100110",
   "11110111001110110110100110100010100000010000101110011111101011111001001110",
   "11110111101110111010011101110000010010100001100100001111110110010010001110",
   "11111000001110111110010101011110001100100001110011100110000000110110011101",
   "11111000101111000010001101101100001110010010011100111001011100101101010010",
   "11111001001111000110000110011010010111110100100000100001011101111111011101",
   "11111001101111001001111111101000101001001000111110110101011011110111001111",
   "11111010001111001101111001010111000010010000111000001100110000100000010101",
   "11111010101111010001110011100101100011001101001100111110111001000111111011",
   "11111011001111010101101110010100001011111110111101100011010101111100101001",
   "11111011101111011001101001100010111100100111001010010001101010001110100110",
   "11111100001111011101100101010001110101000110110011100001011100001111011010",
   "11111100101111100001100001100000110101011110111001101010010101010010000111",
   "11111101001111100101011110001111111101110000011101000100000001101011010001",
   "11111101101111101001011011011111001101111100011110000110010000110000111010",
   "11111110001111101101011001001110100110000011111101001000110100111010100100",
   "11111110101111110001010111011110000110000111111010100011100011100001001110",
   "11111111001111110101010110001101101110001001010110101110010100111111011001",
   "11111111101111111001010101011101011110001001010010000001000100110001000101",
      others => (others => '0'));
      	begin 
      return tmp;
      end init_rom;
	signal rom : memory_t := init_rom;
   signal Y0 :  std_logic_vector(73 downto 0);
begin
	process(clk)
   begin
   if(rising_edge(clk)) then
   	Y0 <= rom(  TO_INTEGER(unsigned(X))  );
   end if;
   end process;
    Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_83_f400_uid128
--                     (IntAdderClassical_83_f400_uid130)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_83_f400_uid128 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(82 downto 0);
          Y : in  std_logic_vector(82 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(82 downto 0)   );
end entity;

architecture arch of IntAdder_83_f400_uid128 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                              LogTable_2_11_66
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity LogTable_2_11_66 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          Y : out  std_logic_vector(65 downto 0)   );
end entity;

architecture arch of LogTable_2_11_66 is
   -- Build a 2-D array type for the RoM
   subtype word_t is std_logic_vector(65 downto 0);
   type memory_t is array(0 to 2047) of word_t;
   function init_rom
      return memory_t is 
      variable tmp : memory_t := (
   "000000000000000000000000000000000000000000000000000100000000000000",
   "000000000010000000000000000000000000000011111000000100000000000000",
   "000000000100000000000000000000000000001111110000000100000000000001",
   "000000000110000000000000000000000000100011101000000100000000000100",
   "000000001000000000000000000000000000111111100000000100000000001011",
   "000000001010000000000000000000000001100011011000000100000000010101",
   "000000001100000000000000000000000010001111010000000100000000100100",
   "000000001110000000000000000000000011000011001000000100000000111001",
   "000000010000000000000000000000000011111111000000000100000001010101",
   "000000010010000000000000000000000101000010111000000100000001111001",
   "000000010100000000000000000000000110001110110000000100000010100110",
   "000000010110000000000000000000000111100010101000000100000011011101",
   "000000011000000000000000000000001000111110100000000100000100011111",
   "000000011010000000000000000000001010100010011000000100000101101101",
   "000000011100000000000000000000001100001110010000000100000111001000",
   "000000011110000000000000000000001110000010001000000100001000110001",
   "000000100000000000000000000000001111111110000000000100001010101001",
   "000000100010000000000000000000010010000001111000000100001100110001",
   "000000100100000000000000000000010100001101110000000100001111001001",
   "000000100110000000000000000000010110100001101000000100010001110100",
   "000000101000000000000000000000011000111101100000000100010100110010",
   "000000101010000000000000000000011011100001011000000100011000000100",
   "000000101100000000000000000000011110001101010000000100011011101011",
   "000000101110000000000000000000100001000001001000000100011111101000",
   "000000110000000000000000000000100011111101000000000100100011111100",
   "000000110010000000000000000000100111000000111000000100101000100111",
   "000000110100000000000000000000101010001100110000000100101101101100",
   "000000110110000000000000000000101101100000101000000100110011001011",
   "000000111000000000000000000000110000111100100000000100111001000101",
   "000000111010000000000000000000110100100000011000000100111111011010",
   "000000111100000000000000000000111000001100010000000101000110001101",
   "000000111110000000000000000000111100000000001000000101001101011110",
   "000001000000000000000000000000111111111100000000000101010101001101",
   "000001000010000000000000000001000011111111111000000101011101011101",
   "000001000100000000000000000001001000001011110000000101100110001110",
   "000001000110000000000000000001001100011111101000000101101111100000",
   "000001001000000000000000000001010000111011100000000101111001010110",
   "000001001010000000000000000001010101011111011000000110000011101111",
   "000001001100000000000000000001011010001011010000000110001110101110",
   "000001001110000000000000000001011110111111001000000110011010010011",
   "000001010000000000000000000001100011111011000000000110100110011110",
   "000001010010000000000000000001101000111110111000000110110011010010",
   "000001010100000000000000000001101110001010110000000111000000101110",
   "000001010110000000000000000001110011011110101000000111001110110101",
   "000001011000000000000000000001111000111010100000000111011101100110",
   "000001011010000000000000000001111110011110011000000111101101000100",
   "000001011100000000000000000010000100001010010000000111111101001110",
   "000001011110000000000000000010001001111110001000001000001110000111",
   "000001100000000000000000000010001111111010000000001000011111101110",
   "000001100010000000000000000010010101111101111000001000110010000101",
   "000001100100000000000000000010011100001001110000001001000101001110",
   "000001100110000000000000000010100010011101101000001001011001001000",
   "000001101000000000000000000010101000111001100000001001101101110110",
   "000001101010000000000000000010101111011101011000001010000011010111",
   "000001101100000000000000000010110110001001010000001010011001101101",
   "000001101110000000000000000010111100111101001000001010110000111010",
   "000001110000000000000000000011000011111001000000001011001000111101",
   "000001110010000000000000000011001010111100111000001011100001111000",
   "000001110100000000000000000011010010001000110000001011111011101100",
   "000001110110000000000000000011011001011100101000001100010110011011",
   "000001111000000000000000000011100000111000100000001100110010000100",
   "000001111010000000000000000011101000011100011000001101001110101001",
   "000001111100000000000000000011110000001000010000001101101100001011",
   "000001111110000000000000000011110111111100001000001110001010101100",
   "000010000000000000000000000011111111111000000000001110101010001011",
   "000010000010000000000000000100000111111011111000001111001010101010",
   "000010000100000000000000000100010000000111110000001111101100001010",
   "000010000110000000000000000100011000011011101000010000001110101100",
   "000010001000000000000000000100100000110111100000010000110010010001",
   "000010001010000000000000000100101001011011011000010001010110111010",
   "000010001100000000000000000100110010000111010000010001111100101000",
   "000010001110000000000000000100111010111011001000010010100011011100",
   "000010010000000000000000000101000011110111000000010011001011011000",
   "000010010010000000000000000101001100111010111000010011110100011011",
   "000010010100000000000000000101010110000110110000010100011110100111",
   "000010010110000000000000000101011111011010101000010101001001111101",
   "000010011000000000000000000101101000110110100000010101110110011110",
   "000010011010000000000000000101110010011010011000010110100100001011",
   "000010011100000000000000000101111100000110010000010111010011000100",
   "000010011110000000000000000110000101111010001000011000000011001100",
   "000010100000000000000000000110001111110110000000011000110100100011",
   "000010100010000000000000000110011001111001111000011001100111001010",
   "000010100100000000000000000110100100000101110000011010011011000010",
   "000010100110000000000000000110101110011001101000011011010000001100",
   "000010101000000000000000000110111000110101100000011100000110101001",
   "000010101010000000000000000111000011011001011000011100111110011010",
   "000010101100000000000000000111001110000101010000011101110111100000",
   "000010101110000000000000000111011000111001001000011110110001111011",
   "000010110000000000000000000111100011110101000000011111101101101110",
   "000010110010000000000000000111101110111000111000100000101010111001",
   "000010110100000000000000000111111010000100110000100001101001011101",
   "000010110110000000000000001000000101011000101000100010101001011010",
   "000010111000000000000000001000010000110100100000100011101010110011",
   "000010111010000000000000001000011100011000011000100100101101101000",
   "000010111100000000000000001000101000000100010000100101110001111010",
   "000010111110000000000000001000110011111000001000100110110111101001",
   "000011000000000000000000001000111111110100000000100111111110111000",
   "000011000010000000000000001001001011110111111000101001000111100111",
   "000011000100000000000000001001011000000011110000101010010001110110",
   "000011000110000000000000001001100100010111101000101011011101101000",
   "000011001000000000000000001001110000110011100000101100101010111101",
   "000011001010000000000000001001111101010111011000101101111001110101",
   "000011001100000000000000001010001010000011010000101111001010010011",
   "000011001110000000000000001010010110110111001000110000011100010110",
   "000011010000000000000000001010100011110011000000110001110000000001",
   "000011010010000000000000001010110000110110111000110011000101010011",
   "000011010100000000000000001010111110000010110000110100011100001111",
   "000011010110000000000000001011001011010110101000110101110100110100",
   "000011011000000000000000001011011000110010100000110111001111000101",
   "000011011010000000000000001011100110010110011000111000101011000001",
   "000011011100000000000000001011110100000010010000111010001000101011",
   "000011011110000000000000001100000001110110001000111011101000000010",
   "000011100000000000000000001100001111110010000000111101001001001001",
   "000011100010000000000000001100011101110101111000111110101011111111",
   "000011100100000000000000001100101100000001110001000000010000100111",
   "000011100110000000000000001100111010010101101001000001110111000000",
   "000011101000000000000000001101001000110001100001000011011111001100",
   "000011101010000000000000001101010111010101011001000101001001001101",
   "000011101100000000000000001101100110000001010001000110110101000010",
   "000011101110000000000000001101110100110101001001001000100010101101",
   "000011110000000000000000001110000011110001000001001010010010010000",
   "000011110010000000000000001110010010110100111001001100000011101010",
   "000011110100000000000000001110100010000000110001001101110110111101",
   "000011110110000000000000001110110001010100101001001111101100001010",
   "000011111000000000000000001111000000110000100001010001100011010011",
   "000011111010000000000000001111010000010100011001010011011100010111",
   "000011111100000000000000001111100000000000010001010101010111011000",
   "000011111110000000000000001111101111110100001001010111010100010111",
   "000100000000000000000000001111111111110000000001011001010011010110",
   "000100000010000000000000010000001111110011111001011011010100010100",
   "000100000100000000000000010000011111111111110001011101010111010011",
   "000100000110000000000000010000110000010011101001011111011100010100",
   "000100001000000000000000010001000000101111100001100001100011011000",
   "000100001010000000000000010001010001010011011001100011101100100000",
   "000100001100000000000000010001100001111111010001100101110111101101",
   "000100001110000000000000010001110010110011001001101000000101000000",
   "000100010000000000000000010010000011101111000001101010010100011010",
   "000100010010000000000000010010010100110010111001101100100101111100",
   "000100010100000000000000010010100101111110110001101110111001100111",
   "000100010110000000000000010010110111010010101001110001001111011100",
   "000100011000000000000000010011001000101110100001110011100111011100",
   "000100011010000000000000010011011010010010011001110110000001101000",
   "000100011100000000000000010011101011111110010001111000011110000001",
   "000100011110000000000000010011111101110010001001111010111100101000",
   "000100100000000000000000010100001111101110000001111101011101011110",
   "000100100010000000000000010100100001110001111010000000000000100100",
   "000100100100000000000000010100110011111101110010000010100101111011",
   "000100100110000000000000010101000110010001101010000101001101100100",
   "000100101000000000000000010101011000101101100010000111110111100000",
   "000100101010000000000000010101101011010001011010001010100011110000",
   "000100101100000000000000010101111101111101010010001101010010010100",
   "000100101110000000000000010110010000110001001010010000000011001111",
   "000100110000000000000000010110100011101101000010010010110110100001",
   "000100110010000000000000010110110110110000111010010101101100001011",
   "000100110100000000000000010111001001111100110010011000100100001110",
   "000100110110000000000000010111011101010000101010011011011110101010",
   "000100111000000000000000010111110000101100100010011110011011100010",
   "000100111010000000000000011000000100010000011010100001011010110110",
   "000100111100000000000000011000010111111100010010100100011100100111",
   "000100111110000000000000011000101011110000001010100111100000110101",
   "000101000000000000000000011000111111101100000010101010100111100011",
   "000101000010000000000000011001010011101111111010101101110000110001",
   "000101000100000000000000011001100111111011110010110000111100011111",
   "000101000110000000000000011001111100001111101010110100001010110000",
   "000101001000000000000000011010010000101011100010110111011011100100",
   "000101001010000000000000011010100101001111011010111010101110111011",
   "000101001100000000000000011010111001111011010010111110000100111000",
   "000101001110000000000000011011001110101111001011000001011101011010",
   "000101010000000000000000011011100011101011000011000100111000100100",
   "000101010010000000000000011011111000101110111011001000010110010101",
   "000101010100000000000000011100001101111010110011001011110110110000",
   "000101010110000000000000011100100011001110101011001111011001110100",
   "000101011000000000000000011100111000101010100011010010111111100100",
   "000101011010000000000000011101001110001110011011010110101000000000",
   "000101011100000000000000011101100011111010010011011010010011001000",
   "000101011110000000000000011101111001101110001011011110000000111110",
   "000101100000000000000000011110001111101010000011100001110001100100",
   "000101100010000000000000011110100101101101111011100101100100111001",
   "000101100100000000000000011110111011111001110011101001011011000000",
   "000101100110000000000000011111010010001101101011101101010011111000",
   "000101101000000000000000011111101000101001100011110001001111100011",
   "000101101010000000000000011111111111001101011011110101001110000011",
   "000101101100000000000000100000010101111001010011111001001111010111",
   "000101101110000000000000100000101100101101001011111101010011100001",
   "000101110000000000000000100001000011101001000100000001011010100011",
   "000101110010000000000000100001011010101100111100000101100100011100",
   "000101110100000000000000100001110001111000110100001001110001001110",
   "000101110110000000000000100010001001001100101100001110000000111011",
   "000101111000000000000000100010100000101000100100010010010011100010",
   "000101111010000000000000100010111000001100011100010110101001000101",
   "000101111100000000000000100011001111111000010100011011000001100101",
   "000101111110000000000000100011100111101100001100011111011101000100",
   "000110000000000000000000100011111111101000000100100011111011100001",
   "000110000010000000000000100100010111101011111100101000011100111110",
   "000110000100000000000000100100101111110111110100101101000001011100",
   "000110000110000000000000100101001000001011101100110001101000111100",
   "000110001000000000000000100101100000100111100100110110010011011111",
   "000110001010000000000000100101111001001011011100111011000001000110",
   "000110001100000000000000100110010001110111010100111111110001110010",
   "000110001110000000000000100110101010101011001101000100100101100100",
   "000110010000000000000000100111000011100111000101001001011100011110",
   "000110010010000000000000100111011100101010111101001110010110011111",
   "000110010100000000000000100111110101110110110101010011010011101001",
   "000110010110000000000000101000001111001010101101011000010011111101",
   "000110011000000000000000101000101000100110100101011101010111011100",
   "000110011010000000000000101001000010001010011101100010011110000111",
   "000110011100000000000000101001011011110110010101100111100111111111",
   "000110011110000000000000101001110101101010001101101100110101000101",
   "000110100000000000000000101010001111100110000101110010000101011010",
   "000110100010000000000000101010101001101001111101110111011000111110",
   "000110100100000000000000101011000011110101110101111100101111110100",
   "000110100110000000000000101011011110001001101110000010001001111100",
   "000110101000000000000000101011111000100101100110000111100111010111",
   "000110101010000000000000101100010011001001011110001101001000000110",
   "000110101100000000000000101100101101110101010110010010101100001010",
   "000110101110000000000000101101001000101001001110011000010011100100",
   "000110110000000000000000101101100011100101000110011101111110010100",
   "000110110010000000000000101101111110101000111110100011101100011101",
   "000110110100000000000000101110011001110100110110101001011101111111",
   "000110110110000000000000101110110101001000101110101111010010111011",
   "000110111000000000000000101111010000100100100110110101001011010010",
   "000110111010000000000000101111101100001000011110111011000111000100",
   "000110111100000000000000110000000111110100010111000001000110010100",
   "000110111110000000000000110000100011101000001111000111001001000010",
   "000111000000000000000000110000111111100100000111001101001111001110",
   "000111000010000000000000110001011011100111111111010011011000111011",
   "000111000100000000000000110001110111110011110111011001100110001001",
   "000111000110000000000000110010010100000111101111011111110110111000",
   "000111001000000000000000110010110000100011100111100110001011001011",
   "000111001010000000000000110011001101000111011111101100100011000010",
   "000111001100000000000000110011101001110011010111110010111110011101",
   "000111001110000000000000110100000110100111001111111001011101011111",
   "000111010000000000000000110100100011100011001000000000000000001000",
   "000111010010000000000000110101000000100111000000000110100110011000",
   "000111010100000000000000110101011101110010111000001101010000010010",
   "000111010110000000000000110101111011000110110000010011111101110101",
   "000111011000000000000000110110011000100010101000011010101111000100",
   "000111011010000000000000110110110110000110100000100001100011111110",
   "000111011100000000000000110111010011110010011000101000011100100110",
   "000111011110000000000000110111110001100110010000101111011000111011",
   "000111100000000000000000111000001111100010001000110110011001000000",
   "000111100010000000000000111000101101100110000000111101011100110100",
   "000111100100000000000000111001001011110001111001000100100100011001",
   "000111100110000000000000111001101010000101110001001011101111110001",
   "000111101000000000000000111010001000100001101001010010111110111011",
   "000111101010000000000000111010100111000101100001011010010001111010",
   "000111101100000000000000111011000101110001011001100001101000101101",
   "000111101110000000000000111011100100100101010001101001000011010110",
   "000111110000000000000000111100000011100001001001110000100001110111",
   "000111110010000000000000111100100010100101000001111000000100001111",
   "000111110100000000000000111101000001110000111001111111101010100000",
   "000111110110000000000000111101100001000100110010000111010100101100",
   "000111111000000000000000111110000000100000101010001111000010110010",
   "000111111010000000000000111110100000000100100010010110110100110100",
   "000111111100000000000000111110111111110000011010011110101010110011",
   "000111111110000000000000111111011111100100010010100110100100110000",
   "001000000000000000000000111111111111100000001010101110100010101101",
   "001000000010000000000001000000011111100100000010110110100100101001",
   "001000000100000000000001000000111111101111111010111110101010100110",
   "001000000110000000000001000001100000000011110011000110110100100101",
   "001000001000000000000001000010000000011111101011001111000010100111",
   "001000001010000000000001000010100001000011100011010111010100101110",
   "001000001100000000000001000011000001101111011011011111101010111000",
   "001000001110000000000001000011100010100011010011101000000101001010",
   "001000010000000000000001000100000011011111001011110000100011100010",
   "001000010010000000000001000100100100100011000011111001000110000010",
   "001000010100000000000001000101000101101110111100000001101100101011",
   "001000010110000000000001000101100111000010110100001010010111011110",
   "001000011000000000000001000110001000011110101100010011000110011100",
   "001000011010000000000001000110101010000010100100011011111001100110",
   "001000011100000000000001000111001011101110011100100100110000111101",
   "001000011110000000000001000111101101100010010100101101101100100010",
   "001000100000000000000001001000001111011110001100110110101100010110",
   "001000100010000000000001001000110001100010000100111111110000011010",
   "001000100100000000000001001001010011101101111101001000111000101111",
   "001000100110000000000001001001110110000001110101010010000101010110",
   "001000101000000000000001001010011000011101101101011011010110010000",
   "001000101010000000000001001010111011000001100101100100101011011110",
   "001000101100000000000001001011011101101101011101101110000101000000",
   "001000101110000000000001001100000000100001010101110111100010111001",
   "001000110000000000000001001100100011011101001110000001000101001001",
   "001000110010000000000001001101000110100001000110001010101011110001",
   "001000110100000000000001001101101001101100111110010100010110110010",
   "001000110110000000000001001110001101000000110110011110000110001100",
   "001000111000000000000001001110110000011100101110100111111010000010",
   "001000111010000000000001001111010100000000100110110001110010010100",
   "001000111100000000000001001111110111101100011110111011101111000011",
   "001000111110000000000001010000011011100000010111000101110000010000",
   "001001000000000000000001010000111111011100001111001111110101111011",
   "001001000010000000000001010001100011100000000111011010000000000111",
   "001001000100000000000001010010000111101011111111100100001110110100",
   "001001000110000000000001010010101011111111110111101110100010000010",
   "001001001000000000000001010011010000011011101111111000111001110100",
   "001001001010000000000001010011110100111111101000000011010110001010",
   "001001001100000000000001010100011001101011100000001101110111000100",
   "001001001110000000000001010100111110011111011000011000011100100101",
   "001001010000000000000001010101100011011011010000100011000110101100",
   "001001010010000000000001010110001000011111001000101101110101011100",
   "001001010100000000000001010110101101101011000000111000101000110100",
   "001001010110000000000001010111010010111110111001000011100000110111",
   "001001011000000000000001010111111000011010110001001110011101100101",
   "001001011010000000000001011000011101111110101001011001011110111110",
   "001001011100000000000001011001000011101010100001100100100101000101",
   "001001011110000000000001011001101001011110011001101111101111111001",
   "001001100000000000000001011010001111011010010001111010111111011101",
   "001001100010000000000001011010110101011110001010000110010011110000",
   "001001100100000000000001011011011011101010000010010001101100110100",
   "001001100110000000000001011100000001111101111010011101001010101011",
   "001001101000000000000001011100101000011001110010101000101101010100",
   "001001101010000000000001011101001110111101101010110100010100110010",
   "001001101100000000000001011101110101101001100011000000000001000100",
   "001001101110000000000001011110011100011101011011001011110010001100",
   "001001110000000000000001011111000011011001010011010111101000001100",
   "001001110010000000000001011111101010011101001011100011100011000011",
   "001001110100000000000001100000010001101001000011101111100010110100",
   "001001110110000000000001100000111000111100111011111011100111011110",
   "001001111000000000000001100001100000011000110100000111110001000011",
   "001001111010000000000001100010000111111100101100010011111111100100",
   "001001111100000000000001100010101111101000100100100000010011000011",
   "001001111110000000000001100011010111011100011100101100101011011111",
   "001010000000000000000001100011111111011000010100111001001000111010",
   "001010000010000000000001100100100111011100001101000101101011010110",
   "001010000100000000000001100101001111101000000101010010010010110010",
   "001010000110000000000001100101110111111011111101011110111111010000",
   "001010001000000000000001100110100000010111110101101011110000110001",
   "001010001010000000000001100111001000111011101101111000100111010110",
   "001010001100000000000001100111110001100111100110000101100011000000",
   "001010001110000000000001101000011010011011011110010010100011110000",
   "001010010000000000000001101001000011010111010110011111101001101000",
   "001010010010000000000001101001101100011011001110101100110100100111",
   "001010010100000000000001101010010101100111000110111010000100101111",
   "001010010110000000000001101010111110111010111111000111011010000001",
   "001010011000000000000001101011101000010110110111010100110100011110",
   "001010011010000000000001101100010001111010101111100010010100000111",
   "001010011100000000000001101100111011100110100111101111111000111101",
   "001010011110000000000001101101100101011010011111111101100011000001",
   "001010100000000000000001101110001111010110011000001011010010010100",
   "001010100010000000000001101110111001011010010000011001000110110111",
   "001010100100000000000001101111100011100110001000100111000000101011",
   "001010100110000000000001110000001101111010000000110100111111110001",
   "001010101000000000000001110000111000010101111001000011000100001010",
   "001010101010000000000001110001100010111001110001010001001101110111",
   "001010101100000000000001110010001101100101101001011111011100111001",
   "001010101110000000000001110010111000011001100001101101110001010000",
   "001010110000000000000001110011100011010101011001111100001011000000",
   "001010110010000000000001110100001110011001010010001010101010000110",
   "001010110100000000000001110100111001100101001010011001001110100110",
   "001010110110000000000001110101100100111001000010100111111000100000",
   "001010111000000000000001110110010000010100111010110110100111110101",
   "001010111010000000000001110110111011111000110011000101011100100110",
   "001010111100000000000001110111100111100100101011010100010110110011",
   "001010111110000000000001111000010011011000100011100011010110011111",
   "001011000000000000000001111000111111010100011011110010011011101010",
   "001011000010000000000001111001101011011000010100000001100110010100",
   "001011000100000000000001111010010111100100001100010000110110100000",
   "001011000110000000000001111011000011111000000100100000001100001110",
   "001011001000000000000001111011110000010011111100101111100111011111",
   "001011001010000000000001111100011100110111110100111111001000010100",
   "001011001100000000000001111101001001100011101101001110101110101101",
   "001011001110000000000001111101110110010111100101011110011010101101",
   "001011010000000000000001111110100011010011011101101110001100010011",
   "001011010010000000000001111111010000010111010101111110000011100010",
   "001011010100000000000001111111111101100011001110001110000000011010",
   "001011010110000000000010000000101010110111000110011110000010111011",
   "001011011000000000000010000001011000010010111110101110001011001000",
   "001011011010000000000010000010000101110110110110111110011001000000",
   "001011011100000000000010000010110011100010101111001110101100100110",
   "001011011110000000000010000011100001010110100111011111000101111010",
   "001011100000000000000010000100001111010010011111101111100100111100",
   "001011100010000000000010000100111101010110011000000000001001101110",
   "001011100100000000000010000101101011100010010000010000110100010010",
   "001011100110000000000010000110011001110110001000100001100100101000",
   "001011101000000000000010000111001000010010000000110010011010110000",
   "001011101010000000000010000111110110110101111001000011010110101100",
   "001011101100000000000010001000100101100001110001010100011000011110",
   "001011101110000000000010001001010100010101101001100101100000000101",
   "001011110000000000000010001010000011010001100001110110101101100100",
   "001011110010000000000010001010110010010101011010001000000000111010",
   "001011110100000000000010001011100001100001010010011001011010001001",
   "001011110110000000000010001100010000110101001010101010111001010010",
   "001011111000000000000010001101000000010001000010111100011110010111",
   "001011111010000000000010001101101111110100111011001110001001010111",
   "001011111100000000000010001110011111100000110011011111111010010100",
   "001011111110000000000010001111001111010100101011110001110001010000",
   "001100000000000000000010001111111111010000100100000011101110001010",
   "001100000010000000000010010000101111010100011100010101110001000100",
   "001100000100000000000010010001011111100000010100100111111010000000",
   "001100000110000000000010010010001111110100001100111010001000111101",
   "001100001000000000000010010011000000010000000101001100011101111101",
   "001100001010000000000010010011110000110011111101011110111001000001",
   "001100001100000000000010010100100001011111110101110001011010001010",
   "001100001110000000000010010101010010010011101110000100000001011010",
   "001100010000000000000010010110000011001111100110010110101110110000",
   "001100010010000000000010010110110100010011011110101001100010001110",
   "001100010100000000000010010111100101011111010110111100011011110101",
   "001100010110000000000010011000010110110011001111001111011011100110",
   "001100011000000000000010011001001000001111000111100010100001100010",
   "001100011010000000000010011001111001110010111111110101101101101010",
   "001100011100000000000010011010101011011110111000001001000000000000",
   "001100011110000000000010011011011101010010110000011100011000100010",
   "001100100000000000000010011100001111001110101000101111110111010101",
   "001100100010000000000010011101000001010010100001000011011100010111",
   "001100100100000000000010011101110011011110011001010111000111101010",
   "001100100110000000000010011110100101110010010001101010111001001111",
   "001100101000000000000010011111011000001110001001111110110001000111",
   "001100101010000000000010100000001010110010000010010010101111010011",
   "001100101100000000000010100000111101011101111010100110110011110100",
   "001100101110000000000010100001110000010001110010111010111110101010",
   "001100110000000000000010100010100011001101101011001111001111111000",
   "001100110010000000000010100011010110010001100011100011100111011110",
   "001100110100000000000010100100001001011101011011111000000101011101",
   "001100110110000000000010100100111100110001010100001100101001110110",
   "001100111000000000000010100101110000001101001100100001010100101010",
   "001100111010000000000010100110100011110001000100110110000101111010",
   "001100111100000000000010100111010111011100111101001010111101100111",
   "001100111110000000000010101000001011010000110101011111111011110010",
   "001101000000000000000010101000111111001100101101110101000000011011",
   "001101000010000000000010101001110011010000100110001010001011100101",
   "001101000100000000000010101010100111011100011110011111011101010000",
   "001101000110000000000010101011011011110000010110110100110101011101",
   "001101001000000000000010101100010000001100001111001010010100001100",
   "001101001010000000000010101101000100110000000111011111111001100000",
   "001101001100000000000010101101111001011011111111110101100101011001",
   "001101001110000000000010101110101110001111111000001011010111111000",
   "001101010000000000000010101111100011001011110000100001010000111101",
   "001101010010000000000010110000011000001111101000110111010000101011",
   "001101010100000000000010110001001101011011100001001101010111000010",
   "001101010110000000000010110010000010101111011001100011100100000010",
   "001101011000000000000010110010111000001011010001111001110111101110",
   "001101011010000000000010110011101101101111001010010000010010000110",
   "001101011100000000000010110100100011011011000010100110110011001010",
   "001101011110000000000010110101011001001110111010111101011010111101",
   "001101100000000000000010110110001111001010110011010100001001011110",
   "001101100010000000000010110111000101001110101011101010111110110000",
   "001101100100000000000010110111111011011010100100000001111010110010",
   "001101100110000000000010111000110001101110011100011000111101100111",
   "001101101000000000000010111001101000001010010100110000000111001110",
   "001101101010000000000010111010011110101110001101000111010111101010",
   "001101101100000000000010111011010101011010000101011110101110111010",
   "001101101110000000000010111100001100001101111101110110001101000001",
   "001101110000000000000010111101000011001001110110001101110001111110",
   "001101110010000000000010111101111010001101101110100101011101110100",
   "001101110100000000000010111110110001011001100110111101010000100010",
   "001101110110000000000010111111101000101101011111010101001010001010",
   "001101111000000000000011000000100000001001010111101101001010101110",
   "001101111010000000000011000001010111101101010000000101010010001110",
   "001101111100000000000011000010001111011001001000011101100000101010",
   "001101111110000000000011000011000111001101000000110101110110000100",
   "001110000000000000000011000011111111001000111001001110010010011110",
   "001110000010000000000011000100110111001100110001100110110101110111",
   "001110000100000000000011000101101111011000101001111111100000010001",
   "001110000110000000000011000110100111101100100010011000010001101110",
   "001110001000000000000011000111100000001000011010110001001010001101",
   "001110001010000000000011001000011000101100010011001010001001110000",
   "001110001100000000000011001001010001011000001011100011010000011000",
   "001110001110000000000011001010001010001100000011111100011110000110",
   "001110010000000000000011001011000011000111111100010101110010111100",
   "001110010010000000000011001011111100001011110100101111001110111001",
   "001110010100000000000011001100110101010111101101001000110001111111",
   "001110010110000000000011001101101110101011100101100010011100001111",
   "001110011000000000000011001110101000000111011101111100001101101010",
   "001110011010000000000011001111100001101011010110010110000110010010",
   "001110011100000000000011010000011011010111001110110000000110000110",
   "001110011110000000000011010001010101001011000111001010001101001000",
   "001110100000000000000011010010001111000110111111100100011011011001",
   "001110100010000000000011010011001001001010110111111110110000111010",
   "001110100100000000000011010100000011010110110000011001001101101100",
   "001110100110000000000011010100111101101010101000110011110001110000",
   "001110101000000000000011010101111000000110100001001110011101000111",
   "001110101010000000000011010110110010101010011001101001001111110010",
   "001110101100000000000011010111101101010110010010000100001001110010",
   "001110101110000000000011011000101000001010001010011111001011001000",
   "001110110000000000000011011001100011000110000010111010010011110101",
   "001110110010000000000011011010011110001001111011010101100011111010",
   "001110110100000000000011011011011001010101110011110000111011011000",
   "001110110110000000000011011100010100101001101100001100011010010000",
   "001110111000000000000011011101010000000101100100101000000000100011",
   "001110111010000000000011011110001011101001011101000011101110010010",
   "001110111100000000000011011111000111010101010101011111100011011110",
   "001110111110000000000011100000000011001001001101111011100000001000",
   "001111000000000000000011100000111111000101000110010111100100010001",
   "001111000010000000000011100001111011001000111110110011101111111010",
   "001111000100000000000011100010110111010100110111010000000011000100",
   "001111000110000000000011100011110011101000101111101100011101101111",
   "001111001000000000000011100100110000000100101000001000111111111110",
   "001111001010000000000011100101101100101000100000100101101001110001",
   "001111001100000000000011100110101001010100011001000010011011001001",
   "001111001110000000000011100111100110001000010001011111010100000110",
   "001111010000000000000011101000100011000100001001111100010100101011",
   "001111010010000000000011101001100000001000000010011001011100111000",
   "001111010100000000000011101010011101010011111010110110101100101110",
   "001111010110000000000011101011011010100111110011010100000100001110",
   "001111011000000000000011101100011000000011101011110001100011011000",
   "001111011010000000000011101101010101100111100100001111001010001111",
   "001111011100000000000011101110010011010011011100101100111000110010",
   "001111011110000000000011101111010001000111010101001010101111000100",
   "001111100000000000000011110000001111000011001101101000101101000101",
   "001111100010000000000011110001001101000111000110000110110010110110",
   "001111100100000000000011110010001011010010111110100101000000010111",
   "001111100110000000000011110011001001100110110111000011010101101011",
   "001111101000000000000011110100001000000010101111100001110010110001",
   "001111101010000000000011110101000110100110101000000000010111101100",
   "001111101100000000000011110110000101010010100000011111000100011100",
   "001111101110000000000011110111000100000110011000111101111001000001",
   "001111110000000000000011111000000011000010010001011100110101011110",
   "001111110010000000000011111001000010000110001001111011111001110010",
   "001111110100000000000011111010000001010010000010011011000110000000",
   "001111110110000000000011111011000000100101111010111010011010000111",
   "001111111000000000000011111100000000000001110011011001110110001010",
   "001111111010000000000011111100111111100101101011111001011010001000",
   "001111111100000000000011111101111111010001100100011001000110000100",
   "001111111110000000000011111110111111000101011100111000111001111101",
   "010000000000000000000011111111111111000001010101011000110101110110",
   "010000000010000000000100000000111111000101001101111000111001101110",
   "010000000100000000000100000001111111010001000110011001000101100111",
   "010000000110000000000100000010111111100100111110111001011001100010",
   "010000001000000000000100000100000000000000110111011001110101100001",
   "010000001010000000000100000101000000100100101111111010011001100100",
   "010000001100000000000100000110000001010000101000011011000101101010",
   "010000001110000000000100000111000010000100100000111011111001111000",
   "010000010000000000000100001000000011000000011001011100110110001100",
   "010000010010000000000100001001000100000100010001111101111010101000",
   "010000010100000000000100001010000101010000001010011111000111001110",
   "010000010110000000000100001011000110100100000011000000011011111101",
   "010000011000000000000100001100000111111111111011100001111000111000",
   "010000011010000000000100001101001001100011110100000011011101111110",
   "010000011100000000000100001110001011001111101100100101001011010001",
   "010000011110000000000100001111001101000011100101000111000000110010",
   "010000100000000000000100010000001110111111011101101000111110100010",
   "010000100010000000000100010001010001000011010110001011000100100010",
   "010000100100000000000100010010010011001111001110101101010010110100",
   "010000100110000000000100010011010101100011000111001111101001010111",
   "010000101000000000000100010100010111111110111111110010001000001101",
   "010000101010000000000100010101011010100010111000010100101111010111",
   "010000101100000000000100010110011101001110110000110111011110110110",
   "010000101110000000000100010111100000000010101001011010010110101011",
   "010000110000000000000100011000100010111110100001111101010110111000",
   "010000110010000000000100011001100110000010011010100000011111011100",
   "010000110100000000000100011010101001001110010011000011110000011000",
   "010000110110000000000100011011101100100010001011100111001001110000",
   "010000111000000000000100011100101111111110000100001010101011100010",
   "010000111010000000000100011101110011100001111100101110010101110000",
   "010000111100000000000100011110110111001101110101010010001000011010",
   "010000111110000000000100011111111011000001101101110110000011100100",
   "010001000000000000000100100000111110111101100110011010000111001100",
   "010001000010000000000100100010000011000001011110111110010011010100",
   "010001000100000000000100100011000111001101010111100010100111111100",
   "010001000110000000000100100100001011100001010000000111000101001000",
   "010001001000000000000100100101001111111101001000101011101010110110",
   "010001001010000000000100100110010100100001000001010000011001000111",
   "010001001100000000000100100111011001001100111001110101001111111110",
   "010001001110000000000100101000011110000000110010011010001111011011",
   "010001010000000000000100101001100010111100101010111111010111011111",
   "010001010010000000000100101010101000000000100011100100101000001010",
   "010001010100000000000100101011101101001100011100001010000001100000",
   "010001010110000000000100101100110010100000010100101111100011011110",
   "010001011000000000000100101101110111111100001101010101001110001000",
   "010001011010000000000100101110111101100000000101111011000001011110",
   "010001011100000000000100110000000011001011111110100000111101100000",
   "010001011110000000000100110001001000111111110111000111000010010010",
   "010001100000000000000100110010001110111011101111101101001111110001",
   "010001100010000000000100110011010100111111101000010011100110000001",
   "010001100100000000000100110100011011001011100000111010000101000010",
   "010001100110000000000100110101100001011111011001100000101100110100",
   "010001101000000000000100110110100111111011010010000111011101011010",
   "010001101010000000000100110111101110011111001010101110010110110100",
   "010001101100000000000100111000110101001011000011010101011001000010",
   "010001101110000000000100111001111011111110111011111100100100000111",
   "010001110000000000000100111011000010111010110100100011111000000010",
   "010001110010000000000100111100001001111110101101001011010100110110",
   "010001110100000000000100111101010001001010100101110010111010100011",
   "010001110110000000000100111110011000011110011110011010101001001010",
   "010001111000000000000100111111011111111010010111000010100000101011",
   "010001111010000000000101000000100111011110001111101010100001001000",
   "010001111100000000000101000001101111001010001000010010101010100011",
   "010001111110000000000101000010110110111110000000111010111100111100",
   "010010000000000000000101000011111110111001111001100011011000010100",
   "010010000010000000000101000101000110111101110010001011111100101011",
   "010010000100000000000101000110001111001001101010110100101010000100",
   "010010000110000000000101000111010111011101100011011101100000011110",
   "010010001000000000000101001000011111111001011100000110011111111100",
   "010010001010000000000101001001101000011101010100101111101000011101",
   "010010001100000000000101001010110001001001001101011000111010000011",
   "010010001110000000000101001011111001111101000110000010010100110000",
   "010010010000000000000101001101000010111000111110101011111000100011",
   "010010010010000000000101001110001011111100110111010101100101011110",
   "010010010100000000000101001111010101001000101111111111011011100011",
   "010010010110000000000101010000011110011100101000101001011010110001",
   "010010011000000000000101010001100111111000100001010011100011001010",
   "010010011010000000000101010010110001011100011001111101110100110000",
   "010010011100000000000101010011111011001000010010101000001111100010",
   "010010011110000000000101010101000100111100001011010010110011100010",
   "010010100000000000000101010110001110111000000011111101100000110010",
   "010010100010000000000101010111011000111011111100101000010111010001",
   "010010100100000000000101011000100011000111110101010011010111000010",
   "010010100110000000000101011001101101011011101101111110100000000100",
   "010010101000000000000101011010110111110111100110101001110010011001",
   "010010101010000000000101011100000010011011011111010101001110000010",
   "010010101100000000000101011101001101000111011000000000110011000000",
   "010010101110000000000101011110010111111011010000101100100001010100",
   "010010110000000000000101011111100010110111001001011000011001000000",
   "010010110010000000000101100000101101111011000010000100011010000011",
   "010010110100000000000101100001111001000110111010110000100100100000",
   "010010110110000000000101100011000100011010110011011100111000010110",
   "010010111000000000000101100100001111110110101100001001010101100110",
   "010010111010000000000101100101011011011010100100110101111100010100",
   "010010111100000000000101100110100111000110011101100010101100011110",
   "010010111110000000000101100111110010111010010110001111100110000110",
   "010011000000000000000101101000111110110110001110111100101001001101",
   "010011000010000000000101101010001010111010000111101001110101110100",
   "010011000100000000000101101011010111000110000000010111001011111100",
   "010011000110000000000101101100100011011001111001000100101011100110",
   "010011001000000000000101101101101111110101110001110010010100110100",
   "010011001010000000000101101110111100011001101010100000000111100100",
   "010011001100000000000101110000001001000101100011001110000011111010",
   "010011001110000000000101110001010101111001011011111100001001110110",
   "010011010000000000000101110010100010110101010100101010011001011010",
   "010011010010000000000101110011101111111001001101011000110010100100",
   "010011010100000000000101110100111101000101000110000111010101011000",
   "010011010110000000000101110110001010011000111110110110000001110110",
   "010011011000000000000101110111010111110100110111100100110111111111",
   "010011011010000000000101111000100101011000110000010011110111110100",
   "010011011100000000000101111001110011000100101001000011000001010110",
   "010011011110000000000101111011000000111000100001110010010100100110",
   "010011100000000000000101111100001110110100011010100001110001100100",
   "010011100010000000000101111101011100111000010011010001011000010100",
   "010011100100000000000101111110101011000100001100000001001000110100",
   "010011100110000000000101111111111001011000000100110001000011000101",
   "010011101000000000000110000001000111110011111101100001000111001010",
   "010011101010000000000110000010010110010111110110010001010101000011",
   "010011101100000000000110000011100101000011101111000001101100110000",
   "010011101110000000000110000100110011110111100111110010001110010100",
   "010011110000000000000110000110000010110011100000100010111001101111",
   "010011110010000000000110000111010001110111011001010011101111000010",
   "010011110100000000000110001000100001000011010010000100101110001110",
   "010011110110000000000110001001110000010111001010110101110111010100",
   "010011111000000000000110001010111111110011000011100111001010010100",
   "010011111010000000000110001100001111010110111100011000100111010001",
   "010011111100000000000110001101011111000010110101001010001110001010",
   "010011111110000000000110001110101110110110101101111011111111000010",
   "010100000000000000000110001111111110110010100110101101111001111001",
   "010100000010000000000110010001001110110110011111011111111110110000",
   "010100000100000000000110010010011111000010011000010010001101100111",
   "010100000110000000000110010011101111010110010001000100100110100001",
   "010100001000000000000110010100111111110010001001110111001001011110",
   "010100001010000000000110010110010000010110000010101001110110011110",
   "010100001100000000000110010111100001000001111011011100101101100100",
   "010100001110000000000110011000110001110101110100001111101110101111",
   "010100010000000000000110011010000010110001101101000010111010000010",
   "010100010010000000000110011011010011110101100101110110001111011100",
   "010100010100000000000110011100100101000001011110101001101111000000",
   "010100010110000000000110011101110110010101010111011101011000101110",
   "010100011000000000000110011111000111110001010000010001001100100110",
   "010100011010000000000110100000011001010101001001000101001010101010",
   "010100011100000000000110100001101011000001000001111001010010111100",
   "010100011110000000000110100010111100110100111010101101100101011011",
   "010100100000000000000110100100001110110000110011100010000010001010",
   "010100100010000000000110100101100000110100101100010110101001001000",
   "010100100100000000000110100110110011000000100101001011011010011000",
   "010100100110000000000110101000000101010100011110000000010101111001",
   "010100101000000000000110101001010111110000010110110101011011101110",
   "010100101010000000000110101010101010010100001111101010101011110110",
   "010100101100000000000110101011111101000000001000100000000110010011",
   "010100101110000000000110101101001111110100000001010101101011000110",
   "010100110000000000000110101110100010101111111010001011011010010001",
   "010100110010000000000110101111110101110011110011000001010011110011",
   "010100110100000000000110110001001000111111101011110111010111101110",
   "010100110110000000000110110010011100010011100100101101100110000100",
   "010100111000000000000110110011101111101111011101100011111110110100",
   "010100111010000000000110110101000011010011010110011010100010000000",
   "010100111100000000000110110110010110111111001111010001001111101010",
   "010100111110000000000110110111101010110011001000001000000111110001",
   "010101000000000000000110111000111110101111000000111111001010010111",
   "010101000010000000000110111010010010110010111001110110010111011110",
   "010101000100000000000110111011100110111110110010101101101111000100",
   "010101000110000000000110111100111011010010101011100101010001001110",
   "010101001000000000000110111110001111101110100100011100111101111010",
   "010101001010000000000110111111100100010010011101010100110101001010",
   "010101001100000000000111000000111000111110010110001100110110111111",
   "010101001110000000000111000010001101110010001111000101000011011010",
   "010101010000000000000111000011100010101110000111111101011010011100",
   "010101010010000000000111000100110111110010000000110101111100000110",
   "010101010100000000000111000110001100111101111001101110101000011010",
   "010101010110000000000111000111100010010001110010100111011111010111",
   "010101011000000000000111001000110111101101101011100000100000111111",
   "010101011010000000000111001010001101010001100100011001101101010011",
   "010101011100000000000111001011100010111101011101010011000100010100",
   "010101011110000000000111001100111000110001010110001100100110000011",
   "010101100000000000000111001110001110101101001111000110010010100001",
   "010101100010000000000111001111100100110001001000000000001001101111",
   "010101100100000000000111010000111010111101000000111010001011101110",
   "010101100110000000000111010010010001010000111001110100011000011111",
   "010101101000000000000111010011100111101100110010101110110000000011",
   "010101101010000000000111010100111110010000101011101001010010011011",
   "010101101100000000000111010110010100111100100100100011111111101000",
   "010101101110000000000111010111101011110000011101011110110111101011",
   "010101110000000000000111011001000010101100010110011001111010100101",
   "010101110010000000000111011010011001110000001111010101001000010111",
   "010101110100000000000111011011110000111100001000010000100001000010",
   "010101110110000000000111011101001000010000000001001100000100100110",
   "010101111000000000000111011110011111101011111010000111110011000110",
   "010101111010000000000111011111110111001111110011000011101100100010",
   "010101111100000000000111100001001110111011101011111111110000111011",
   "010101111110000000000111100010100110101111100100111100000000010010",
   "010110000000000000000111100011111110101011011101111000011010101000",
   "010110000010000000000111100101010110101111010110110100111111111110",
   "010110000100000000000111100110101110111011001111110001110000010100",
   "010110000110000000000111101000000111001111001000101110101011101101",
   "010110001000000000000111101001011111101011000001101011110010001001",
   "010110001010000000000111101010111000001110111010101001000011101000",
   "010110001100000000000111101100010000111010110011100110100000001110",
   "010110001110000000000111101101101001101110101100100100000111111000",
   "010110010000000000000111101111000010101010100101100001111010101010",
   "010110010010000000000111110000011011101110011110011111111000100100",
   "010110010100000000000111110001110100111010010111011110000001100110",
   "010110010110000000000111110011001110001110010000011100010101110011",
   "010110011000000000000111110100100111101010001001011010110101001010",
   "010110011010000000000111110110000001001110000010011001011111101110",
   "010110011100000000000111110111011010111001111011011000010101011111",
   "010110011110000000000111111000110100101101110100010111010110011110",
   "010110100000000000000111111010001110101001101101010110100010101011",
   "010110100010000000000111111011101000101101100110010101111010001001",
   "010110100100000000000111111101000010111001011111010101011100111000",
   "010110100110000000000111111110011101001101011000010101001010111000",
   "010110101000000000000111111111110111101001010001010101000100001100",
   "010110101010000000001000000001010010001101001010010101001000110011",
   "010110101100000000001000000010101100111001000011010101011000110000",
   "010110101110000000001000000100000111101100111100010101110100000010",
   "010110110000000000001000000101100010101000110101010110011010101100",
   "010110110010000000001000000110111101101100101110010111001100101101",
   "010110110100000000001000001000011000111000100111011000001010001000",
   "010110110110000000001000001001110100001100100000011001010010111100",
   "010110111000000000001000001011001111101000011001011010100111001100",
   "010110111010000000001000001100101011001100010010011100000110110111",
   "010110111100000000001000001110000110111000001011011101110010000000",
   "010110111110000000001000001111100010101100000100011111101000100110",
   "010111000000000000001000010000111110100111111101100001101010101100",
   "010111000010000000001000010010011010101011110110100011111000010001",
   "010111000100000000001000010011110110110111101111100110010001010111",
   "010111000110000000001000010101010011001011101000101000110110000000",
   "010111001000000000001000010110101111100111100001101011100110001011",
   "010111001010000000001000011000001100001011011010101110100001111010",
   "010111001100000000001000011001101000110111010011110001101001001110",
   "010111001110000000001000011011000101101011001100110100111100001001",
   "010111010000000000001000011100100010100111000101111000011010101010",
   "010111010010000000001000011101111111101010111110111100000100110100",
   "010111010100000000001000011111011100110110110111111111111010100110",
   "010111010110000000001000100000111010001010110001000011111100000010",
   "010111011000000000001000100010010111100110101010001000001001001010",
   "010111011010000000001000100011110101001010100011001100100001111100",
   "010111011100000000001000100101010010110110011100010001000110011101",
   "010111011110000000001000100110110000101010010101010101110110101011",
   "010111100000000000001000101000001110100110001110011010110010101000",
   "010111100010000000001000101001101100101010000111011111111010010110",
   "010111100100000000001000101011001010110110000000100101001101110100",
   "010111100110000000001000101100101001001001111001101010101101000100",
   "010111101000000000001000101110000111100101110010110000011000000111",
   "010111101010000000001000101111100110001001101011110110001110111110",
   "010111101100000000001000110001000100110101100100111100010001101010",
   "010111101110000000001000110010100011101001011110000010100000001100",
   "010111110000000000001000110100000010100101010111001000111010100110",
   "010111110010000000001000110101100001101001010000001111100000110110",
   "010111110100000000001000110111000000110101001001010110010011000001",
   "010111110110000000001000111000100000001001000010011101010001000101",
   "010111111000000000001000111001111111100100111011100100011011000100",
   "010111111010000000001000111011011111001000110100101011110000111111",
   "010111111100000000001000111100111110110100101101110011010010110111",
   "010111111110000000001000111110011110101000100110111011000000101101",
   "011000000000000000001000111111111110100100100000000010111010100010",
   "011000000010000000001001000001011110101000011001001011000000010111",
   "011000000100000000001001000010111110110100010010010011010010001101",
   "011000000110000000001001000100011111001000001011011011110000000101",
   "011000001000000000001001000101111111100100000100100100011010000000",
   "011000001010000000001001000111100000000111111101101101001111111111",
   "011000001100000000001001001001000000110011110110110110010010000011",
   "011000001110000000001001001010100001100111101111111111100000001101",
   "011000010000000000001001001100000010100011101001001000111010011110",
   "011000010010000000001001001101100011100111100010010010100000110110",
   "011000010100000000001001001111000100110011011011011100010011011000",
   "011000010110000000001001010000100110000111010100100110010010000100",
   "011000011000000000001001010010000111100011001101110000011100111100",
   "011000011010000000001001010011101001000111000110111010110011111110",
   "011000011100000000001001010101001010110011000000000101010111001110",
   "011000011110000000001001010110101100100110111001010000000110101100",
   "011000100000000000001001011000001110100010110010011011000010011000",
   "011000100010000000001001011001110000100110101011100110001010010110",
   "011000100100000000001001011011010010110010100100110001011110100100",
   "011000100110000000001001011100110101000110011101111100111111000011",
   "011000101000000000001001011110010111100010010111001000101011110110",
   "011000101010000000001001011111111010000110010000010100100100111100",
   "011000101100000000001001100001011100110010001001100000101010011000",
   "011000101110000000001001100010111111100110000010101100111100001010",
   "011000110000000000001001100100100010100001111011111001011010010011",
   "011000110010000000001001100110000101100101110101000110000100110100",
   "011000110100000000001001100111101000110001101110010010111011101101",
   "011000110110000000001001101001001100000101100111011111111111000001",
   "011000111000000000001001101010101111100001100000101101001110110000",
   "011000111010000000001001101100010011000101011001111010101010111010",
   "011000111100000000001001101101110110110001010011001000010011100010",
   "011000111110000000001001101111011010100101001100010110001000101000",
   "011001000000000000001001110000111110100001000101100100001010001100",
   "011001000010000000001001110010100010100100111110110010011000010001",
   "011001000100000000001001110100000110110000111000000000110010110110",
   "011001000110000000001001110101101011000100110001001111011001111110",
   "011001001000000000001001110111001111100000101010011110001101101000",
   "011001001010000000001001111000110100000100100011101101001101110111",
   "011001001100000000001001111010011000110000011100111100011010101010",
   "011001001110000000001001111011111101100100010110001011110100000100",
   "011001010000000000001001111101100010100000001111011011011010000100",
   "011001010010000000001001111111000111100100001000101011001100101101",
   "011001010100000000001010000000101100110000000001111011001011111111",
   "011001010110000000001010000010010010000011111011001011010111111010",
   "011001011000000000001010000011110111011111110100011011110000100000",
   "011001011010000000001010000101011101000011101101101100010101110011",
   "011001011100000000001010000111000010101111100110111101000111110010",
   "011001011110000000001010001000101000100011100000001110000110100000",
   "011001100000000000001010001010001110011111011001011111010001111100",
   "011001100010000000001010001011110100100011010010110000101010001001",
   "011001100100000000001010001101011010101111001100000010001111000110",
   "011001100110000000001010001111000001000011000101010100000000110110",
   "011001101000000000001010010000100111011110111110100101111111011000",
   "011001101010000000001010010010001110000010110111111000001010101110",
   "011001101100000000001010010011110100101110110001001010100010111010",
   "011001101110000000001010010101011011100010101010011101000111111100",
   "011001110000000000001010010111000010011110100011101111111001110100",
   "011001110010000000001010011000101001100010011101000010111000100100",
   "011001110100000000001010011010010000101110010110010110000100001101",
   "011001110110000000001010011011111000000010001111101001011100110000",
   "011001111000000000001010011101011111011110001000111101000010001111",
   "011001111010000000001010011111000111000010000010010000110100101001",
   "011001111100000000001010100000101110101101111011100100110100000000",
   "011001111110000000001010100010010110100001110100111001000000010110",
   "011010000000000000001010100011111110011101101110001101011001101010",
   "011010000010000000001010100101100110100001100111100001111111111110",
   "011010000100000000001010100111001110101101100000110110110011010100",
   "011010000110000000001010101000110111000001011010001011110011101010",
   "011010001000000000001010101010011111011101010011100001000001000100",
   "011010001010000000001010101100001000000001001100110110011011100011",
   "011010001100000000001010101101110000101101000110001100000011000110",
   "011010001110000000001010101111011001100000111111100001110111110000",
   "011010010000000000001010110001000010011100111000110111111001100000",
   "011010010010000000001010110010101011100000110010001110001000011000",
   "011010010100000000001010110100010100101100101011100100100100011000",
   "011010010110000000001010110101111110000000100100111011001101100100",
   "011010011000000000001010110111100111011100011110010010000011111010",
   "011010011010000000001010111001010001000000010111101001000111011100",
   "011010011100000000001010111010111010101100010001000000011000001011",
   "011010011110000000001010111100100100100000001010010111110110001000",
   "011010100000000000001010111110001110011100000011101111100001010100",
   "011010100010000000001010111111111000011111111101000111011001110000",
   "011010100100000000001011000001100010101011110110011111011111011110",
   "011010100110000000001011000011001100111111101111110111110010011100",
   "011010101000000000001011000100110111011011101001010000010010101110",
   "011010101010000000001011000110100001111111100010101001000000010100",
   "011010101100000000001011001000001100101011011100000001111011010000",
   "011010101110000000001011001001110111011111010101011011000011100000",
   "011010110000000000001011001011100010011011001110110100011001001000",
   "011010110010000000001011001101001101011111001000001101111100001000",
   "011010110100000000001011001110111000101011000001100111101100100001",
   "011010110110000000001011010000100011111110111011000001101010010100",
   "011010111000000000001011010010001111011010110100011011110101100010",
   "011010111010000000001011010011111010111110101101110110001110001100",
   "011010111100000000001011010101100110101010100111010000110100010011",
   "011010111110000000001011010111010010011110100000101011100111111000",
   "011011000000000000001011011000111110011010011010000110101000111100",
   "011011000010000000001011011010101010011110010011100001110111100000",
   "011011000100000000001011011100010110101010001100111101010011100100",
   "011011000110000000001011011110000010111110000110011000111101001011",
   "011011001000000000001011011111101111011001111111110100110100010101",
   "011011001010000000001011100001011011111101111001010000111001000011",
   "011011001100000000001011100011001000101001110010101101001011010110",
   "011011001110000000001011100100110101011101101100001001101011001110",
   "011011010000000000001011100110100010011001100101100110011000101110",
   "011011010010000000001011101000001111011101011111000011010011110110",
   "011011010100000000001011101001111100101001011000100000011100100110",
   "011011010110000000001011101011101001111101010001111101110011000010",
   "011011011000000000001011101101010111011001001011011011010111000111",
   "011011011010000000001011101111000100111101000100111001001000111001",
   "011011011100000000001011110000110010101000111110010111001000011000",
   "011011011110000000001011110010100000011100110111110101010101100100",
   "011011100000000000001011110100001110011000110001010011110000100000",
   "011011100010000000001011110101111100011100101010110010011001001100",
   "011011100100000000001011110111101010101000100100010001001111101000",
   "011011100110000000001011111001011000111100011101110000010011110111",
   "011011101000000000001011111011000111011000010111001111100101111000",
   "011011101010000000001011111100110101111100010000101111000101101110",
   "011011101100000000001011111110100100101000001010001110110011011001",
   "011011101110000000001100000000010011011100000011101110101110111010",
   "011011110000000000001100000010000010010111111101001110111000010001",
   "011011110010000000001100000011110001011011110110101111001111100000",
   "011011110100000000001100000101100000100111110000001111110100101010",
   "011011110110000000001100000111001111111011101001110000100111101100",
   "011011111000000000001100001000111111010111100011010001101000101010",
   "011011111010000000001100001010101110111011011100110010110111100011",
   "011011111100000000001100001100011110100111010110010100010100011010",
   "011011111110000000001100001110001110011011001111110101111111001110",
   "011100000000000000001100001111111110010111001001010111111000000010",
   "011100000010000000001100010001101110011011000010111001111110110101",
   "011100000100000000001100010011011110100110111100011100010011101010",
   "011100000110000000001100010101001110111010110101111110110110100000",
   "011100001000000000001100010110111111010110101111100001100111011010",
   "011100001010000000001100011000101111111010101001000100100110010111",
   "011100001100000000001100011010100000100110100010100111110011011010",
   "011100001110000000001100011100010001011010011100001011001110100010",
   "011100010000000000001100011110000010010110010101101110110111110001",
   "011100010010000000001100011111110011011010001111010010101111001000",
   "011100010100000000001100100001100100100110001000110110110100101001",
   "011100010110000000001100100011010101111010000010011011001000010100",
   "011100011000000000001100100101000111010101111011111111101010001001",
   "011100011010000000001100100110111000111001110101100100011010001010",
   "011100011100000000001100101000101010100101101111001001011000011000",
   "011100011110000000001100101010011100011001101000101110100100110101",
   "011100100000000000001100101100001110010101100010010011111111100000",
   "011100100010000000001100101110000000011001011011111001101000011100",
   "011100100100000000001100101111110010100101010101011111011111101000",
   "011100100110000000001100110001100100111001001111000101100101000110",
   "011100101000000000001100110011010111010101001000101011111000111000",
   "011100101010000000001100110101001001111001000010010010011010111100",
   "011100101100000000001100110110111100100100111011111001001011010111",
   "011100101110000000001100111000101111011000110101100000001010001000",
   "011100110000000000001100111010100010010100101111000111010111001110",
   "011100110010000000001100111100010101011000101000101110110010101110",
   "011100110100000000001100111110001000100100100010010110011100100110",
   "011100110110000000001100111111111011111000011011111110010100111000",
   "011100111000000000001101000001101111010100010101100110011011100110",
   "011100111010000000001101000011100010111000001111001110110000101110",
   "011100111100000000001101000101010110100100001000110111010100010101",
   "011100111110000000001101000111001010011000000010100000000110011001",
   "011101000000000000001101001000111110010011111100001001000110111100",
   "011101000010000000001101001010110010010111110101110010010110000000",
   "011101000100000000001101001100100110100011101111011011110011100100",
   "011101000110000000001101001110011010110111101001000101011111101010",
   "011101001000000000001101010000001111010011100010101111011010010010",
   "011101001010000000001101010010000011110111011100011001100011100000",
   "011101001100000000001101010011111000100011010110000011111011010010",
   "011101001110000000001101010101101101010111001111101110100001101010",
   "011101010000000000001101010111100010010011001001011001010110101001",
   "011101010010000000001101011001010111010111000011000100011010010000",
   "011101010100000000001101011011001100100010111100101111101100100000",
   "011101010110000000001101011101000001110110110110011011001101011010",
   "011101011000000000001101011110110111010010110000000110111100111111",
   "011101011010000000001101100000101100110110101001110010111011010000",
   "011101011100000000001101100010100010100010100011011111001000001110",
   "011101011110000000001101100100011000010110011101001011100011111010",
   "011101100000000000001101100110001110010010010110111000001110010101",
   "011101100010000000001101101000000100010110010000100101000111100000",
   "011101100100000000001101101001111010100010001010010010001111011100",
   "011101100110000000001101101011110000110110000011111111100110001010",
   "011101101000000000001101101101100111010001111101101101001011101011",
   "011101101010000000001101101111011101110101110111011011000000000000",
   "011101101100000000001101110001010100100001110001001001000011001010",
   "011101101110000000001101110011001011010101101010110111010101001010",
   "011101110000000000001101110101000010010001100100100101110110000000",
   "011101110010000000001101110110111001010101011110010100100101110000",
   "011101110100000000001101111000110000100001011000000011100100011000",
   "011101110110000000001101111010100111110101010001110010110001111010",
   "011101111000000000001101111100011111010001001011100010001110010110",
   "011101111010000000001101111110010110110101000101010001111001101111",
   "011101111100000000001110000000001110100000111111000001110100000101",
   "011101111110000000001110000010000110010100111000110001111101011001",
   "011110000000000000001110000011111110010000110010100010010101101100",
   "011110000010000000001110000101110110010100101100010010111100111110",
   "011110000100000000001110000111101110100000100110000011110011010010",
   "011110000110000000001110001001100110110100011111110100111000101000",
   "011110001000000000001110001011011111010000011001100110001101000001",
   "011110001010000000001110001101010111110100010011010111110000011110",
   "011110001100000000001110001111010000100000001101001001100011000000",
   "011110001110000000001110010001001001010100000110111011100100100111",
   "011110010000000000001110010011000010010000000000101101110101010110",
   "011110010010000000001110010100111011010011111010100000010101001100",
   "011110010100000000001110010110110100011111110100010011000100001100",
   "011110010110000000001110011000101101110011101110000110000010010110",
   "011110011000000000001110011010100111001111100111111001001111101010",
   "011110011010000000001110011100100000110011100001101100101100001100",
   "011110011100000000001110011110011010011111011011100000010111111001",
   "011110011110000000001110100000010100010011010101010100010010110100",
   "011110100000000000001110100010001110001111001111001000011101000000",
   "011110100010000000001110100100001000010011001000111100110110011010",
   "011110100100000000001110100110000010011111000010110001011111000110",
   "011110100110000000001110100111111100110010111100100110010111000011",
   "011110101000000000001110101001110111001110110110011011011110010100",
   "011110101010000000001110101011110001110010110000010000110100111000",
   "011110101100000000001110101101101100011110101010000110011010110010",
   "011110101110000000001110101111100111010010100011111100010000000010",
   "011110110000000000001110110001100010001110011101110010010100101000",
   "011110110010000000001110110011011101010010010111101000101000100110",
   "011110110100000000001110110101011000011110010001011111001011111110",
   "011110110110000000001110110111010011110010001011010101111110110000",
   "011110111000000000001110111001001111001110000101001101000000111100",
   "011110111010000000001110111011001010110001111111000100010010100101",
   "011110111100000000001110111101000110011101111000111011110011101010",
   "011110111110000000001110111111000010010001110010110011100100001110",
   "011111000000000000001111000000111110001101101100101011100100010000",
   "011111000010000000001111000010111010010001100110100011110011110011",
   "011111000100000000001111000100110110011101100000011100010010110110",
   "011111000110000000001111000110110010110001011010010101000001011100",
   "011111001000000000001111001000101111001101010100001101111111100100",
   "011111001010000000001111001010101011110001001110000111001101010000",
   "011111001100000000001111001100101000011101001000000000101010100010",
   "011111001110000000001111001110100101010001000001111010010111011010",
   "011111010000000000001111010000100010001100111011110100010011111000",
   "011111010010000000001111010010011111010000110101101110011111111110",
   "011111010100000000001111010100011100011100101111101000111011101110",
   "011111010110000000001111010110011001110000101001100011100111000111",
   "011111011000000000001111011000010111001100100011011110100010001100",
   "011111011010000000001111011010010100110000011101011001101100111100",
   "011111011100000000001111011100010010011100010111010101000111011001",
   "011111011110000000001111011110010000010000010001010000110001100100",
   "011111100000000000001111100000001110001100001011001100101011011111",
   "011111100010000000001111100010001100010000000101001000110101001001",
   "011111100100000000001111100100001010011011111111000101001110100100",
   "011111100110000000001111100110001000101111111001000001110111110010",
   "011111101000000000001111101000000111001011110010111110110000110010",
   "011111101010000000001111101010000101101111101100111011111001100110",
   "011111101100000000001111101100000100011011100110111001010010010000",
   "011111101110000000001111101110000011001111100000110110111010101111",
   "011111110000000000001111110000000010001011011010110100110011000101",
   "011111110010000000001111110010000001001111010100110010111011010100",
   "011111110100000000001111110100000000011011001110110001010011011010",
   "011111110110000000001111110101111111101111001000101111111011011100",
   "011111111000000000001111110111111111001011000010101110110011011000",
   "011111111010000000001111111001111110101110111100101101111011010000",
   "011111111100000000001111111011111110011010110110101101010011000110",
   "011111111110000000001111111101111110001110110000101100111010111000",
   "100000000000000000001111111111111110001010101010101100110010101011",
   "100000000010000000010000000001111110001110100100101100111010011101",
   "100000000100000000010000000011111110011010011110101101010010010000",
   "100000000110000000010000000101111110101110011000101101111010000101",
   "100000001000000000010000000111111111001010010010101110110001111101",
   "100000001010000000010000001001111111101110001100101111111001111001",
   "100000001100000000010000001100000000011010000110110001010001111011",
   "100000001110000000010000001110000001001110000000110010111010000010",
   "100000010000000000010000010000000010001001111010110100110010010000",
   "100000010010000000010000010010000011001101110100110110111010100110",
   "100000010100000000010000010100000100011001101110111001010011000101",
   "100000010110000000010000010110000101101101101000111011111011101110",
   "100000011000000000010000011000000111001001100010111110110100100010",
   "100000011010000000010000011010001000101101011101000001111101100010",
   "100000011100000000010000011100001010011001010111000101010110101111",
   "100000011110000000010000011110001100001101010001001001000000001010",
   "100000100000000000010000100000001110001001001011001100111001110100",
   "100000100010000000010000100010010000001101000101010001000011101110",
   "100000100100000000010000100100010010011000111111010101011101111001",
   "100000100110000000010000100110010100101100111001011010001000010110",
   "100000101000000000010000101000010111001000110011011111000011000110",
   "100000101010000000010000101010011001101100101101100100001110001010",
   "100000101100000000010000101100011100011000100111101001101001100011",
   "100000101110000000010000101110011111001100100001101111010101010010",
   "100000110000000000010000110000100010001000011011110101010001011000",
   "100000110010000000010000110010100101001100010101111011011101110110",
   "100000110100000000010000110100101000011000010000000001111010101101",
   "100000110110000000010000110110101011101100001010001000100111111110",
   "100000111000000000010000111000101111001000000100001111100101101010",
   "100000111010000000010000111010110010101011111110010110110011110010",
   "100000111100000000010000111100110110010111111000011110010010010110",
   "100000111110000000010000111110111010001011110010100110000001011001",
   "100001000000000000010001000000111110000111101100101110000000111011",
   "100001000010000000010001000011000010001011100110110110010000111101",
   "100001000100000000010001000101000110010111100000111110110001100000",
   "100001000110000000010001000111001010101011011011000111100010100101",
   "100001001000000000010001001001001111000111010101010000100100001101",
   "100001001010000000010001001011010011101011001111011001110110011000",
   "100001001100000000010001001101011000010111001001100011011001001001",
   "100001001110000000010001001111011101001011000011101101001100100000",
   "100001010000000000010001010001100010000110111101110111010000011110",
   "100001010010000000010001010011100111001010111000000001100101000100",
   "100001010100000000010001010101101100010110110010001100001010010010",
   "100001010110000000010001010111110001101010101100010111000000001011",
   "100001011000000000010001011001110111000110100110100010000110101111",
   "100001011010000000010001011011111100101010100000101101011101111111",
   "100001011100000000010001011110000010010110011010111001000101111011",
   "100001011110000000010001100000001000001010010101000100111110100110",
   "100001100000000000010001100010001110000110001111010001001000000000",
   "100001100010000000010001100100010100001010001001011101100010001001",
   "100001100100000000010001100110011010010110000011101010001101000100",
   "100001100110000000010001101000100000101001111101110111001000110001",
   "100001101000000000010001101010100111000101111000000100010101010000",
   "100001101010000000010001101100101101101001110010010001110010100100",
   "100001101100000000010001101110110100010101101100011111100000101101",
   "100001101110000000010001110000111011001001100110101101011111101011",
   "100001110000000000010001110011000010000101100000111011101111100001",
   "100001110010000000010001110101001001001001011011001010010000001111",
   "100001110100000000010001110111010000010101010101011001000001110101",
   "100001110110000000010001111001010111101001001111101000000100010110",
   "100001111000000000010001111011011111000101001001110111010111110010",
   "100001111010000000010001111101100110101001000100000110111100001001",
   "100001111100000000010001111111101110010100111110010110110001011110",
   "100001111110000000010010000001110110001000111000100110110111110000",
   "100010000000000000010010000011111110000100110010110111001111000010",
   "100010000010000000010010000110000110001000101101000111110111010011",
   "100010000100000000010010001000001110010100100111011000110000100110",
   "100010000110000000010010001010010110101000100001101001111010111011",
   "100010001000000000010010001100011111000100011011111011010110010010",
   "100010001010000000010010001110100111101000010110001101000010101110",
   "100010001100000000010010010000110000010100010000011111000000001110",
   "100010001110000000010010010010111001001000001010110001001110110101",
   "100010010000000000010010010101000010000100000101000011101110100010",
   "100010010010000000010010010111001011000111111111010110011111011000",
   "100010010100000000010010011001010100010011111001101001100001010110",
   "100010010110000000010010011011011101100111110011111100110100011111",
   "100010011000000000010010011101100111000011101110010000011000110010",
   "100010011010000000010010011111110000100111101000100100001110010010",
   "100010011100000000010010100001111010010011100010111000010100111110",
   "100010011110000000010010100100000100000111011101001100101100111000",
   "100010100000000000010010100110001110000011010111100001010110000010",
   "100010100010000000010010101000011000000111010001110110010000011011",
   "100010100100000000010010101010100010010011001100001011011100000110",
   "100010100110000000010010101100101100100111000110100000111001000010",
   "100010101000000000010010101110110111000011000000110110100111010001",
   "100010101010000000010010110001000001100110111011001100100110110101",
   "100010101100000000010010110011001100010010110101100010110111101101",
   "100010101110000000010010110101010111000110101111111001011001111100",
   "100010110000000000010010110111100010000010101010010000001101100001",
   "100010110010000000010010111001101101000110100100100111010010011110",
   "100010110100000000010010111011111000010010011110111110101000110101",
   "100010110110000000010010111110000011100110011001010110010000100101",
   "100010111000000000010011000000001111000010010011101110001001110000",
   "100010111010000000010011000010011010100110001110000110010100011000",
   "100010111100000000010011000100100110010010001000011110110000011100",
   "100010111110000000010011000110110010000110000010110111011101111110",
   "100011000000000000010011001000111110000001111101010000011100111111",
   "100011000010000000010011001011001010000101110111101001101101100001",
   "100011000100000000010011001101010110010001110010000011001111100011",
   "100011000110000000010011001111100010100101101100011101000011000111",
   "100011001000000000010011010001101111000001100110110111001000001111",
   "100011001010000000010011010011111011100101100001010001011110111010",
   "100011001100000000010011010110001000010001011011101100000111001010",
   "100011001110000000010011011000010101000101010110000111000001000000",
   "100011010000000000010011011010100010000001010000100010001100011101",
   "100011010010000000010011011100101111000101001010111101101001100011",
   "100011010100000000010011011110111100010001000101011001011000010001",
   "100011010110000000010011100001001001100100111111110101011000101001",
   "100011011000000000010011100011010111000000111010010001101010101100",
   "100011011010000000010011100101100100100100110100101110001110011011",
   "100011011100000000010011100111110010010000101111001011000011111000",
   "100011011110000000010011101010000000000100101001101000001011000010",
   "100011100000000000010011101100001110000000100100000101100011111011",
   "100011100010000000010011101110011100000100011110100011001110100100",
   "100011100100000000010011110000101010010000011001000001001010111110",
   "100011100110000000010011110010111000100100010011011111011001001010",
   "100011101000000000010011110101000111000000001101111101111001001001",
   "100011101010000000010011110111010101100100001000011100101010111101",
   "100011101100000000010011111001100100010000000010111011101110100101",
   "100011101110000000010011111011110011000011111101011011000100000011",
   "100011110000000000010011111110000001111111110111111010101011011000",
   "100011110010000000010100000000010001000011110010011010100100100101",
   "100011110100000000010100000010100000001111101100111010101111101011",
   "100011110110000000010100000100101111100011100111011011001100101011",
   "100011111000000000010100000110111110111111100001111011111011100110",
   "100011111010000000010100001001001110100011011100011100111100011101",
   "100011111100000000010100001011011110001111010110111110001111010001",
   "100011111110000000010100001101101110000011010001011111110100000011",
   "100100000000000000010100001111111101111111001100000001101010110100",
   "100100000010000000010100010010001110000011000110100011110011100101",
   "100100000100000000010100010100011110001111000001000110001110010111",
   "100100000110000000010100010110101110100010111011101000111011001011",
   "100100001000000000010100011000111110111110110110001011111010000010",
   "100100001010000000010100011011001111100010110000101111001010111101",
   "100100001100000000010100011101100000001110101011010010101101111101",
   "100100001110000000010100011111110001000010100101110110100011000011",
   "100100010000000000010100100010000001111110100000011010101010010000",
   "100100010010000000010100100100010011000010011010111111000011100101",
   "100100010100000000010100100110100100001110010101100011101111000011",
   "100100010110000000010100101000110101100010010000001000101100101011",
   "100100011000000000010100101011000110111110001010101101111100011110",
   "100100011010000000010100101101011000100010000101010011011110011101",
   "100100011100000000010100101111101010001101111111111001010010101001",
   "100100011110000000010100110001111100000001111010011111011001000011",
   "100100100000000000010100110100001101111101110101000101110001101011",
   "100100100010000000010100110110100000000001101111101100011100100100",
   "100100100100000000010100111000110010001101101010010011011001101110",
   "100100100110000000010100111011000100100001100100111010101001001010",
   "100100101000000000010100111101010110111101011111100010001010111001",
   "100100101010000000010100111111101001100001011010001001111110111100",
   "100100101100000000010101000001111100001101010100110010000101010100",
   "100100101110000000010101000100001111000001001111011010011110000001",
   "100100110000000000010101000110100001111101001010000011001001000110",
   "100100110010000000010101001000110101000001000100101100000110100011",
   "100100110100000000010101001011001000001100111111010101010110011001",
   "100100110110000000010101001101011011100000111001111110111000101001",
   "100100111000000000010101001111101110111100110100101000101101010011",
   "100100111010000000010101010010000010100000101111010010110100011010",
   "100100111100000000010101010100010110001100101001111101001101111110",
   "100100111110000000010101010110101010000000100100100111111010000000",
   "100101000000000000010101011000111101111100011111010010111000100001",
   "100101000010000000010101011011010010000000011001111110001001100001",
   "100101000100000000010101011101100110001100010100101001101101000011",
   "100101000110000000010101011111111010100000001111010101100011000111",
   "100101001000000000010101100010001110111100001010000001101011101110",
   "100101001010000000010101100100100011100000000100101110000110111000",
   "100101001100000000010101100110111000001011111111011010110100101000",
   "100101001110000000010101101001001100111111111010000111110100111110",
   "100101010000000000010101101011100001111011110100110101000111111010",
   "100101010010000000010101101101110110111111101111100010101101011111",
   "100101010100000000010101110000001100001011101010010000100101101101",
   "100101010110000000010101110010100001011111100100111110110000100100",
   "100101011000000000010101110100110110111011011111101101001110000111",
   "100101011010000000010101110111001100011111011010011011111110010110",
   "100101011100000000010101111001100010001011010101001011000001010001",
   "100101011110000000010101111011110111111111001111111010010110111011",
   "100101100000000000010101111110001101111011001010101001111111010100",
   "100101100010000000010110000000100011111111000101011001111010011100",
   "100101100100000000010110000010111010001011000000001010001000010110",
   "100101100110000000010110000101010000011110111010111010101001000010",
   "100101101000000000010110000111100110111010110101101011011100100000",
   "100101101010000000010110001001111101011110110000011100100010110011",
   "100101101100000000010110001100010100001010101011001101111011111010",
   "100101101110000000010110001110101010111110100101111111100111111000",
   "100101110000000000010110010001000001111010100000110001100110101101",
   "100101110010000000010110010011011000111110011011100011111000011001",
   "100101110100000000010110010101110000001010010110010110011100111111",
   "100101110110000000010110011000000111011110010001001001010100011110",
   "100101111000000000010110011010011110111010001011111100011110111001",
   "100101111010000000010110011100110110011110000110101111111100001111",
   "100101111100000000010110011111001110001010000001100011101100100011",
   "100101111110000000010110100001100101111101111100010111101111110100",
   "100110000000000000010110100011111101111001110111001100000110000101",
   "100110000010000000010110100110010101111101110010000000101111010101",
   "100110000100000000010110101000101110001001101100110101101011100111",
   "100110000110000000010110101011000110011101100111101010111010111010",
   "100110001000000000010110101101011110111001100010100000011101010001",
   "100110001010000000010110101111110111011101011101010110010010101011",
   "100110001100000000010110110010010000001001011000001100011011001011",
   "100110001110000000010110110100101000111101010011000010110110110000",
   "100110010000000000010110110111000001111001001101111001100101011101",
   "100110010010000000010110111001011010111101001000110000100111010001",
   "100110010100000000010110111011110100001001000011100111111100001111",
   "100110010110000000010110111110001101011100111110011111100100010110",
   "100110011000000000010111000000100110111000111001010111011111101001",
   "100110011010000000010111000011000000011100110100001111101110000111",
   "100110011100000000010111000101011010001000101111001000001111110010",
   "100110011110000000010111000111110011111100101010000001000100101100",
   "100110100000000000010111001010001101111000100100111010001100110100",
   "100110100010000000010111001100100111111100011111110011101000001101",
   "100110100100000000010111001111000010001000011010101101010110110110",
   "100110100110000000010111010001011100011100010101100111011000110001",
   "100110101000000000010111010011110110111000010000100001101110000000",
   "100110101010000000010111010110010001011100001011011100010110100010",
   "100110101100000000010111011000101100001000000110010111010010011001",
   "100110101110000000010111011011000110111100000001010010100001100111",
   "100110110000000000010111011101100001110111111100001110000100001011",
   "100110110010000000010111011111111100111011110111001001111010001000",
   "100110110100000000010111100010011000000111110010000110000011011101",
   "100110110110000000010111100100110011011011101101000010100000001100",
   "100110111000000000010111100111001110110111100111111111010000010111",
   "100110111010000000010111101001101010011011100010111100010011111101",
   "100110111100000000010111101100000110000111011101111001101011000000",
   "100110111110000000010111101110100001111011011000110111010101100001",
   "100111000000000000010111110000111101110111010011110101010011100010",
   "100111000010000000010111110011011001111011001110110011100101000010",
   "100111000100000000010111110101110110000111001001110010001010000011",
   "100111000110000000010111111000010010011011000100110001000010100111",
   "100111001000000000010111111010101110110110111111110000001110101101",
   "100111001010000000010111111101001011011010111010101111101110010111",
   "100111001100000000010111111111101000000110110101101111100001100110",
   "100111001110000000011000000010000100111010110000101111101000011100",
   "100111010000000000011000000100100001110110101011110000000010111000",
   "100111010010000000011000000110111110111010100110110000110000111100",
   "100111010100000000011000001001011100000110100001110001110010101001",
   "100111010110000000011000001011111001011010011100110011001000000000",
   "100111011000000000011000001110010110110110010111110100110001000011",
   "100111011010000000011000010000110100011010010010110110101101110001",
   "100111011100000000011000010011010010000110001101111000111110001100",
   "100111011110000000011000010101101111111010001000111011100010010101",
   "100111100000000000011000011000001101110110000011111110011010001101",
   "100111100010000000011000011010101011111001111111000001100101110110",
   "100111100100000000011000011101001010000101111010000101000101001111",
   "100111100110000000011000011111101000011001110101001000111000011010",
   "100111101000000000011000100010000110110101110000001100111111011000",
   "100111101010000000011000100100100101011001101011010001011010001010",
   "100111101100000000011000100111000100000101100110010110001000110001",
   "100111101110000000011000101001100010111001100001011011001011001111",
   "100111110000000000011000101100000001110101011100100000100001100011",
   "100111110010000000011000101110100000111001010111100110001011101111",
   "100111110100000000011000110001000000000101010010101100001001110100",
   "100111110110000000011000110011011111011001001101110010011011110011",
   "100111111000000000011000110101111110110101001000111001000001101101",
   "100111111010000000011000111000011110011001000011111111111011100011",
   "100111111100000000011000111010111110000100111111000111001001010110",
   "100111111110000000011000111101011101111000111010001110101011000111",
   "101000000000000000011000111111111101110100110101010110100000110111",
   "101000000010000000011001000010011101111000110000011110101010101000",
   "101000000100000000011001000100111110000100101011100111001000011001",
   "101000000110000000011001000111011110011000100110101111111010001100",
   "101000001000000000011001001001111110110100100001111001000000000010",
   "101000001010000000011001001100011111011000011101000010011001111100",
   "101000001100000000011001001111000000000100011000001100000111111011",
   "101000001110000000011001010001100000111000010011010110001010000000",
   "101000010000000000011001010100000001110100001110100000100000001100",
   "101000010010000000011001010110100010111000001001101011001010100000",
   "101000010100000000011001011001000100000100000100110110001000111101",
   "101000010110000000011001011011100101011000000000000001011011100100",
   "101000011000000000011001011110000110110011111011001101000010010110",
   "101000011010000000011001100000101000010111110110011000111101010100",
   "101000011100000000011001100011001010000011110001100101001100011111",
   "101000011110000000011001100101101011110111101100110001101111111000",
   "101000100000000000011001101000001101110011100111111110100111100000",
   "101000100010000000011001101010101111110111100011001011110011011000",
   "101000100100000000011001101101010010000011011110011001010011100001",
   "101000100110000000011001101111110100010111011001100111000111111100",
   "101000101000000000011001110010010110110011010100110101010000101010",
   "101000101010000000011001110100111001010111010000000011101101101100",
   "101000101100000000011001110111011100000011001011010010011111000010",
   "101000101110000000011001111001111110110111000110100001100100101111",
   "101000110000000000011001111100100001110011000001110000111110110011",
   "101000110010000000011001111111000100110110111101000000101101001111",
   "101000110100000000011010000001101000000010111000010000110000000100",
   "101000110110000000011010000100001011010110110011100001000111010011",
   "101000111000000000011010000110101110110010101110110001110010111101",
   "101000111010000000011010001001010010010110101010000010110011000011",
   "101000111100000000011010001011110110000010100101010100000111100110",
   "101000111110000000011010001110011001110110100000100101110000100111",
   "101001000000000000011010010000111101110010011011110111101110000111",
   "101001000010000000011010010011100001110110010111001010000000000110",
   "101001000100000000011010010110000110000010010010011100100110100111",
   "101001000110000000011010011000101010010110001101101111100001101010",
   "101001001000000000011010011011001110110010001001000010110001010000",
   "101001001010000000011010011101110011010110000100010110010101011010",
   "101001001100000000011010100000011000000001111111101010001110001001",
   "101001001110000000011010100010111100110101111010111110011011011101",
   "101001010000000000011010100101100001110001110110010010111101011001",
   "101001010010000000011010101000000110110101110001100111110011111101",
   "101001010100000000011010101010101100000001101100111100111111001010",
   "101001010110000000011010101101010001010101101000010010011111000001",
   "101001011000000000011010101111110110110001100011101000010011100011",
   "101001011010000000011010110010011100010101011110111110011100110000",
   "101001011100000000011010110101000010000001011010010100111010101011",
   "101001011110000000011010110111100111110101010101101011101101010100",
   "101001100000000000011010111010001101110001010001000010110100101100",
   "101001100010000000011010111100110011110101001100011010010000110100",
   "101001100100000000011010111111011010000001000111110010000001101100",
   "101001100110000000011011000010000000010101000011001010000111010111",
   "101001101000000000011011000100100110110000111110100010100001110101",
   "101001101010000000011011000111001101010100111001111011010001000111",
   "101001101100000000011011001001110100000000110101010100010101001101",
   "101001101110000000011011001100011010110100110000101101101110001010",
   "101001110000000000011011001111000001110000101100000111011011111110",
   "101001110010000000011011010001101000110100100111100001011110101010",
   "101001110100000000011011010100010000000000100010111011110110001110",
   "101001110110000000011011010110110111010100011110010110100010101101",
   "101001111000000000011011011001011110110000011001110001100100000111",
   "101001111010000000011011011100000110010100010101001100111010011100",
   "101001111100000000011011011110101110000000010000101000100101101111",
   "101001111110000000011011100001010101110100001100000100100110000000",
   "101010000000000000011011100011111101110000000111100000111011001111",
   "101010000010000000011011100110100101110100000010111101100101011111",
   "101010000100000000011011101001001101111111111110011010100100110000",
   "101010000110000000011011101011110110010011111001110111111001000011",
   "101010001000000000011011101110011110101111110101010101100010011000",
   "101010001010000000011011110001000111010011110000110011100000110010",
   "101010001100000000011011110011101111111111101100010001110100010001",
   "101010001110000000011011110110011000110011100111110000011100110101",
   "101010010000000000011011111001000001101111100011001111011010100001",
   "101010010010000000011011111011101010110011011110101110101101010100",
   "101010010100000000011011111110010011111111011010001110010101010001",
   "101010010110000000011100000000111101010011010101101110010010011000",
   "101010011000000000011100000011100110101111010001001110100100101001",
   "101010011010000000011100000110010000010011001100101111001100000111",
   "101010011100000000011100001000111001111111001000010000001000110010",
   "101010011110000000011100001011100011110011000011110001011010101010",
   "101010100000000000011100001110001101101110111111010011000001110010",
   "101010100010000000011100010000110111110010111010110100111110001001",
   "101010100100000000011100010011100001111110110110010111001111110010",
   "101010100110000000011100010110001100010010110001111001110110101101",
   "101010101000000000011100011000110110101110101101011100110010111010",
   "101010101010000000011100011011100001010010101001000000000100011100",
   "101010101100000000011100011110001011111110100100100011101011010010",
   "101010101110000000011100100000110110110010100000000111100111011111",
   "101010110000000000011100100011100001101110011011101011111001000010",
   "101010110010000000011100100110001100110010010111010000011111111110",
   "101010110100000000011100101000110111111110010010110101011100010011",
   "101010110110000000011100101011100011010010001110011010101110000001",
   "101010111000000000011100101110001110101110001010000000010101001011",
   "101010111010000000011100110000111010010010000101100110010001110000",
   "101010111100000000011100110011100101111110000001001100100011110011",
   "101010111110000000011100110110010001110001111100110011001011010011",
   "101011000000000000011100111000111101101101111000011010001000010011",
   "101011000010000000011100111011101001110001110100000001011010110010",
   "101011000100000000011100111110010101111101101111101001000010110011",
   "101011000110000000011101000001000010010001101011010001000000010101",
   "101011001000000000011101000011101110101101100110111001010011011011",
   "101011001010000000011101000110011011010001100010100001111100000100",
   "101011001100000000011101001001000111111101011110001010111010010011",
   "101011001110000000011101001011110100110001011001110100001110000111",
   "101011010000000000011101001110100001101101010101011101110111100011",
   "101011010010000000011101010001001110110001010001000111110110100110",
   "101011010100000000011101010011111011111101001100110010001011010011",
   "101011010110000000011101010110101001010001001000011100110101101001",
   "101011011000000000011101011001010110101101000100000111110101101011",
   "101011011010000000011101011100000100010000111111110011001011011000",
   "101011011100000000011101011110110001111100111011011110110110110011",
   "101011011110000000011101100001011111110000110111001010110111111011",
   "101011100000000000011101100100001101101100110010110111001110110010",
   "101011100010000000011101100110111011110000101110100011111011011010",
   "101011100100000000011101101001101001111100101010010000111101110010",
   "101011100110000000011101101100011000010000100101111110010101111101",
   "101011101000000000011101101111000110101100100001101100000011111010",
   "101011101010000000011101110001110101010000011101011010000111101100",
   "101011101100000000011101110100100011111100011001001000100001010010",
   "101011101110000000011101110111010010110000010100110111010000101110",
   "101011110000000000011101111010000001101100010000100110010110000010",
   "101011110010000000011101111100110000110000001100010101110001001101",
   "101011110100000000011101111111011111111100001000000101100010010010",
   "101011110110000000011110000010001111010000000011110101101001010000",
   "101011111000000000011110000100111110101011111111100110000110001001",
   "101011111010000000011110000111101110001111111011010110111000111111",
   "101011111100000000011110001010011101111011110111001000000001110001",
   "101011111110000000011110001101001101101111110010111001100000100010",
   "101100000000000000011110001111111101101011101110101011010101010001",
   "101100000010000000011110010010101101101111101010011101100000000000",
   "101100000100000000011110010101011101111011100110010000000000110001",
   "101100000110000000011110011000001110001111100010000010110111100011",
   "101100001000000000011110011010111110101011011101110110000100011000",
   "101100001010000000011110011101101111001111011001101001100111010010",
   "101100001100000000011110100000011111111011010101011101100000010000",
   "101100001110000000011110100011010000101111010001010001101111010100",
   "101100010000000000011110100110000001101011001101000110010100100000",
   "101100010010000000011110101000110010101111001000111011001111110011",
   "101100010100000000011110101011100011111011000100110000100001001111",
   "101100010110000000011110101110010101001111000000100110001000110110",
   "101100011000000000011110110001000110101010111100011100000110100111",
   "101100011010000000011110110011111000001110111000010010011010100100",
   "101100011100000000011110110110101001111010110100001001000100101111",
   "101100011110000000011110111001011011101110110000000000000101000111",
   "101100100000000000011110111100001101101010101011110111011011101110",
   "101100100010000000011110111110111111101110100111101111001000100101",
   "101100100100000000011111000001110001111010100011100111001011101110",
   "101100100110000000011111000100100100001110011111011111100101001000",
   "101100101000000000011111000111010110101010011011011000010100110101",
   "101100101010000000011111001010001001001110010111010001011010110111",
   "101100101100000000011111001100111011111010010011001010110111001101",
   "101100101110000000011111001111101110101110001111000100101001111001",
   "101100110000000000011111010010100001101010001010111110110010111100",
   "101100110010000000011111010101010100101110000110111001010010011000",
   "101100110100000000011111011000000111111010000010110100001000001100",
   "101100110110000000011111011010111011001101111110101111010100011010",
   "101100111000000000011111011101101110101001111010101010110111000011",
   "101100111010000000011111100000100010001101110110100110110000001001",
   "101100111100000000011111100011010101111001110010100010111111101011",
   "101100111110000000011111100110001001101101101110011111100101101011",
   "101101000000000000011111101000111101101001101010011100100010001010",
   "101101000010000000011111101011110001101101100110011001110101001010",
   "101101000100000000011111101110100101111001100010010111011110101010",
   "101101000110000000011111110001011010001101011110010101011110101100",
   "101101001000000000011111110100001110101001011010010011110101010001",
   "101101001010000000011111110111000011001101010110010010100010011010",
   "101101001100000000011111111001110111111001010010010001100110001001",
   "101101001110000000011111111100101100101101001110010001000000011101",
   "101101010000000000011111111111100001101001001010010000110001011000",
   "101101010010000000100000000010010110101101000110010000111000111011",
   "101101010100000000100000000101001011111001000010010001010111000111",
   "101101010110000000100000001000000001001100111110010010001011111110",
   "101101011000000000100000001010110110101000111010010011010111011111",
   "101101011010000000100000001101101100001100110110010100111001101100",
   "101101011100000000100000010000100001111000110010010110110010100110",
   "101101011110000000100000010011010111101100101110011001000010001110",
   "101101100000000000100000010110001101101000101010011011101000100110",
   "101101100010000000100000011001000011101100100110011110100101101101",
   "101101100100000000100000011011111001111000100010100001111001100101",
   "101101100110000000100000011110110000001100011110100101100100001111",
   "101101101000000000100000100001100110101000011010101001100101101100",
   "101101101010000000100000100100011101001100010110101101111101111101",
   "101101101100000000100000100111010011111000010010110010101101000011",
   "101101101110000000100000101010001010101100001110110111110011000000",
   "101101110000000000100000101101000001101000001010111101001111110011",
   "101101110010000000100000101111111000101100000111000011000011011110",
   "101101110100000000100000110010101111111000000011001001001110000010",
   "101101110110000000100000110101100111001011111111001111101111100000",
   "101101111000000000100000111000011110100111111011010110100111111001",
   "101101111010000000100000111011010110001011110111011101110111001110",
   "101101111100000000100000111110001101110111110011100101011101100000",
   "101101111110000000100001000001000101101011101111101101011010110001",
   "101110000000000000100001000011111101100111101011110101101111000000",
   "101110000010000000100001000110110101101011100111111110011010001111",
   "101110000100000000100001001001101101110111100100000111011100011111",
   "101110000110000000100001001100100110001011100000010000110101110001",
   "101110001000000000100001001111011110100111011100011010100110000110",
   "101110001010000000100001010010010111001011011000100100101101011111",
   "101110001100000000100001010101001111110111010100101111001011111101",
   "101110001110000000100001011000001000101011010000111010000001100001",
   "101110010000000000100001011011000001100111001101000101001110001100",
   "101110010010000000100001011101111010101011001001010000110010000000",
   "101110010100000000100001100000110011110111000101011100101100111100",
   "101110010110000000100001100011101101001011000001101000111111000010",
   "101110011000000000100001100110100110100110111101110101101000010011",
   "101110011010000000100001101001100000001010111010000010101000110000",
   "101110011100000000100001101100011001110110110110010000000000011010",
   "101110011110000000100001101111010011101010110010011101101111010010",
   "101110100000000000100001110010001101100110101110101011110101011001",
   "101110100010000000100001110101000111101010101010111010010010110000",
   "101110100100000000100001111000000001110110100111001001000111011000",
   "101110100110000000100001111010111100001010100011011000010011010010",
   "101110101000000000100001111101110110100110011111100111110110011111",
   "101110101010000000100010000000110001001010011011110111110001000000",
   "101110101100000000100010000011101011110110011000001000000010110110",
   "101110101110000000100010000110100110101010010100011000101100000010",
   "101110110000000000100010001001100001100110010000101001101100100101",
   "101110110010000000100010001100011100101010001100111011000100100000",
   "101110110100000000100010001111010111110110001001001100110011110100",
   "101110110110000000100010010010010011001010000101011110111010100010",
   "101110111000000000100010010101001110100110000001110001011000101011",
   "101110111010000000100010011000001010001001111110000100001110010000",
   "101110111100000000100010011011000101110101111010010111011011010010",
   "101110111110000000100010011110000001101001110110101010111111110010",
   "101111000000000000100010100000111101100101110010111110111011110001",
   "101111000010000000100010100011111001101001101111010011001111010000",
   "101111000100000000100010100110110101110101101011100111111010010000",
   "101111000110000000100010101001110010001001100111111100111100110010",
   "101111001000000000100010101100101110100101100100010010010110110111",
   "101111001010000000100010101111101011001001100000101000001000100000",
   "101111001100000000100010110010100111110101011100111110010001101110",
   "101111001110000000100010110101100100101001011001010100110010100010",
   "101111010000000000100010111000100001100101010101101011101010111101",
   "101111010010000000100010111011011110101001010010000010111011000000",
   "101111010100000000100010111110011011110101001110011010100010101100",
   "101111010110000000100011000001011001001001001010110010100010000010",
   "101111011000000000100011000100010110100101000111001010111001000011",
   "101111011010000000100011000111010100001001000011100011100111110000",
   "101111011100000000100011001010010001110100111111111100101110001010",
   "101111011110000000100011001101001111101000111100010110001100010010",
   "101111100000000000100011010000001101100100111000110000000010001001",
   "101111100010000000100011010011001011101000110101001010001111110000",
   "101111100100000000100011010110001001110100110001100100110101001000",
   "101111100110000000100011011001001000001000101101111111110010010010",
   "101111101000000000100011011100000110100100101010011011000111001111",
   "101111101010000000100011011111000101001000100110110110110100000000",
   "101111101100000000100011100010000011110100100011010010111000100110",
   "101111101110000000100011100101000010101000011111101111010101000010",
   "101111110000000000100011101000000001100100011100001100001001010101",
   "101111110010000000100011101011000000101000011000101001010101100000",
   "101111110100000000100011101101111111110100010101000110111001100100",
   "101111110110000000100011110000111111001000010001100100110101100001",
   "101111111000000000100011110011111110100100001110000011001001011010",
   "101111111010000000100011110110111110001000001010100001110101001111",
   "101111111100000000100011111001111101110100000111000000111001000001",
   "101111111110000000100011111100111101101000000011100000010100110001",
   "110000000000000000100011111111111101100100000000000000001000100000",
   "110000000010000000100100000010111101100111111100100000010100001111",
   "110000000100000000100100000101111101110011111001000000110111111111",
   "110000000110000000100100001000111110000111110101100001110011110001",
   "110000001000000000100100001011111110100011110010000011000111100110",
   "110000001010000000100100001110111111000111101110100100110011011111",
   "110000001100000000100100010001111111110011101011000110110111011101",
   "110000001110000000100100010101000000100111100111101001010011100000",
   "110000010000000000100100011000000001100011100100001100000111101011",
   "110000010010000000100100011011000010100111100000101111010011111110",
   "110000010100000000100100011110000011110011011101010010111000011010",
   "110000010110000000100100100001000101000111011001110110110101000000",
   "110000011000000000100100100100000110100011010110011011001001110001",
   "110000011010000000100100100111001000000111010010111111110110101110",
   "110000011100000000100100101010001001110011001111100100111011111000",
   "110000011110000000100100101101001011100111001100001010011001010000",
   "110000100000000000100100110000001101100011001000110000001110110110",
   "110000100010000000100100110011001111100111000101010110011100101101",
   "110000100100000000100100110110010001110011000001111101000010110101",
   "110000100110000000100100111001010100000110111110100100000001001111",
   "110000101000000000100100111100010110100010111011001011010111111100",
   "110000101010000000100100111111011001000110110111110011000110111101",
   "110000101100000000100101000010011011110010110100011011001110010011",
   "110000101110000000100101000101011110100110110001000011101101111111",
   "110000110000000000100101001000100001100010101101101100100110000001",
   "110000110010000000100101001011100100100110101010010101110110011100",
   "110000110100000000100101001110100111110010100110111111011111010000",
   "110000110110000000100101010001101011000110100011101001100000011110",
   "110000111000000000100101010100101110100010100000010011111010000111",
   "110000111010000000100101010111110010000110011100111110101100001100",
   "110000111100000000100101011010110101110010011001101001110110101110",
   "110000111110000000100101011101111001100110010110010101011001101101",
   "110001000000000000100101100000111101100010010011000001010101001100",
   "110001000010000000100101100100000001100110001111101101101001001011",
   "110001000100000000100101100111000101110010001100011010010101101011",
   "110001000110000000100101101010001010000110001001000111011010101101",
   "110001001000000000100101101101001110100010000101110100111000010010",
   "110001001010000000100101110000010011000110000010100010101110011010",
   "110001001100000000100101110011010111110001111111010000111101001000",
   "110001001110000000100101110110011100100101111011111111100100011100",
   "110001010000000000100101111001100001100001111000101110100100010111",
   "110001010010000000100101111100100110100101110101011101111100111010",
   "110001010100000000100101111111101011110001110010001101101110000110",
   "110001010110000000100110000010110001000101101110111101110111111011",
   "110001011000000000100110000101110110100001101011101110011010011100",
   "110001011010000000100110001000111100000101101000011111010101101001",
   "110001011100000000100110001100000001110001100101010000101001100011",
   "110001011110000000100110001111000111100101100010000010010110001011",
   "110001100000000000100110010010001101100001011110110100011011100010",
   "110001100010000000100110010101010011100101011011100110111001101000",
   "110001100100000000100110011000011001110001011000011001110000100000",
   "110001100110000000100110011011100000000101010101001101000000001010",
   "110001101000000000100110011110100110100001010010000000101000100111",
   "110001101010000000100110100001101101000101001110110100101001111000",
   "110001101100000000100110100100110011110001001011101001000011111101",
   "110001101110000000100110100111111010100101001000011101110110111001",
   "110001110000000000100110101011000001100001000101010011000010101100",
   "110001110010000000100110101110001000100101000010001000100111010111",
   "110001110100000000100110110001001111110000111110111110100100111011",
   "110001110110000000100110110100010111000100111011110100111011011001",
   "110001111000000000100110110111011110100000111000101011101010110001",
   "110001111010000000100110111010100110000100110101100010110011000110",
   "110001111100000000100110111101101101110000110010011010010100011000",
   "110001111110000000100111000000110101100100101111010010001110101000",
   "110010000000000000100111000011111101100000101100001010100001110111",
   "110010000010000000100111000111000101100100101001000011001110000101",
   "110010000100000000100111001010001101110000100101111100010011010101",
   "110010000110000000100111001101010110000100100010110101110001100111",
   "110010001000000000100111010000011110100000011111101111101000111100",
   "110010001010000000100111010011100111000100011100101001111001010100",
   "110010001100000000100111010110101111110000011001100100100010110010",
   "110010001110000000100111011001111000100100010110011111100101010110",
   "110010010000000000100111011101000001100000010011011011000001000001",
   "110010010010000000100111100000001010100100010000010110110101110100",
   "110010010100000000100111100011010011110000001101010011000011101111",
   "110010010110000000100111100110011101000100001010001111101010110101",
   "110010011000000000100111101001100110100000000111001100101011000110",
   "110010011010000000100111101100110000000100000100001010000100100011",
   "110010011100000000100111101111111001110000000001000111110111001101",
   "110010011110000000100111110011000011100011111110000110000011000100",
   "110010100000000000100111110110001101011111111011000100101000001011",
   "110010100010000000100111111001010111100011111000000011100110100010",
   "110010100100000000100111111100100001101111110101000010111110001010",
   "110010100110000000100111111111101100000011110010000010101111000011",
   "110010101000000000101000000010110110011111101111000010111001010000",
   "110010101010000000101000000110000001000011101100000011011100110001",
   "110010101100000000101000001001001011101111101001000100011001100111",
   "110010101110000000101000001100010110100011100110000101101111110011",
   "110010110000000000101000001111100001011111100011000111011111010101",
   "110010110010000000101000010010101100100011100000001001101000010000",
   "110010110100000000101000010101110111101111011101001100001010100100",
   "110010110110000000101000011001000011000011011010001111000110010010",
   "110010111000000000101000011100001110011111010111010010011011011010",
   "110010111010000000101000011111011010000011010100010110001001111111",
   "110010111100000000101000100010100101101111010001011010010010000001",
   "110010111110000000101000100101110001100011001110011110110011100001",
   "110011000000000000101000101000111101011111001011100011101110011111",
   "110011000010000000101000101100001001100011001000101001000010111110",
   "110011000100000000101000101111010101101111000101101110110000111110",
   "110011000110000000101000110010100010000011000010110100111000100000",
   "110011001000000000101000110101101110011110111111111011011001100100",
   "110011001010000000101000111000111011000010111101000010010100001101",
   "110011001100000000101000111100000111101110111010001001101000011011",
   "110011001110000000101000111111010100100010110111010001010110001111",
   "110011010000000000101001000010100001011110110100011001011101101001",
   "110011010010000000101001000101101110100010110001100001111110101100",
   "110011010100000000101001001000111011101110101110101010111001011000",
   "110011010110000000101001001100001001000010101011110100001101101110",
   "110011011000000000101001001111010110011110101000111101111011101111",
   "110011011010000000101001010010100100000010100110001000000011011011",
   "110011011100000000101001010101110001101110100011010010100100110101",
   "110011011110000000101001011000111111100010100000011101011111111101",
   "110011100000000000101001011100001101011110011101101000110100110100",
   "110011100010000000101001011111011011100010011010110100100011011010",
   "110011100100000000101001100010101001101110011000000000101011110010",
   "110011100110000000101001100101111000000010010101001101001101111100",
   "110011101000000000101001101001000110011110010010011010001001111001",
   "110011101010000000101001101100010101000010001111100111011111101001",
   "110011101100000000101001101111100011101110001100110101001111001111",
   "110011101110000000101001110010110010100010001010000011011000101011",
   "110011110000000000101001110110000001011110000111010001111011111110",
   "110011110010000000101001111001010000100010000100100000111001001000",
   "110011110100000000101001111100011111101110000001110000010000001100",
   "110011110110000000101001111111101111000001111111000000000001001010",
   "110011111000000000101010000010111110011101111100010000001100000011",
   "110011111010000000101010000110001110000001111001100000110000110111",
   "110011111100000000101010001001011101101101110110110001101111101001",
   "110011111110000000101010001100101101100001110100000011001000011001",
   "110100000000000000101010001111111101011101110001010100111011001000",
   "110100000010000000101010010011001101100001101110100111000111110110",
   "110100000100000000101010010110011101101101101011111001101110100110",
   "110100000110000000101010011001101110000001101001001100101111011000",
   "110100001000000000101010011100111110011101100110100000001010001101",
   "110100001010000000101010100000001111000001100011110011111111000101",
   "110100001100000000101010100011011111101101100001001000001110000011",
   "110100001110000000101010100110110000100001011110011100110111000111",
   "110100010000000000101010101010000001011101011011110001111010010010",
   "110100010010000000101010101101010010100001011001000111010111100100",
   "110100010100000000101010110000100011101101010110011101001111000000",
   "110100010110000000101010110011110101000001010011110011100000100110",
   "110100011000000000101010110111000110011101010001001010001100010111",
   "110100011010000000101010111010011000000001001110100001010010010011",
   "110100011100000000101010111101101001101101001011111000110010011101",
   "110100011110000000101011000000111011100001001001010000101100110101",
   "110100100000000000101011000100001101011101000110101001000001011100",
   "110100100010000000101011000111011111100001000100000001110000010010",
   "110100100100000000101011001010110001101101000001011010111001011010",
   "110100100110000000101011001110000100000000111110110100011100110100",
   "110100101000000000101011010001010110011100111100001110011010100001",
   "110100101010000000101011010100101001000000111001101000110010100001",
   "110100101100000000101011010111111011101100110111000011100100110111",
   "110100101110000000101011011011001110100000110100011110110001100011",
   "110100110000000000101011011110100001011100110001111010011000100110",
   "110100110010000000101011100001110100100000101111010110011010000000",
   "110100110100000000101011100101000111101100101100110010110101110100",
   "110100110110000000101011101000011011000000101010001111101100000010",
   "110100111000000000101011101011101110011100100111101100111100101011",
   "110100111010000000101011101111000010000000100101001010100111101111",
   "110100111100000000101011110010010101101100100010101000101101010001",
   "110100111110000000101011110101101001100000100000000111001101010001",
   "110101000000000000101011111000111101011100011101100110000111110000",
   "110101000010000000101011111100010001100000011011000101011100101110",
   "110101000100000000101011111111100101101100011000100101001100001110",
   "110101000110000000101100000010111010000000010110000101010110010000",
   "110101001000000000101100000110001110011100010011100101111010110101",
   "110101001010000000101100001001100011000000010001000110111001111101",
   "110101001100000000101100001100110111101100001110101000010011101011",
   "110101001110000000101100010000001100100000001100001010000111111111",
   "110101010000000000101100010011100001011100001001101100010110111010",
   "110101010010000000101100010110110110100000000111001111000000011100",
   "110101010100000000101100011010001011101100000100110010000100101000",
   "110101010110000000101100011101100001000000000010010101100011011110",
   "110101011000000000101100100000110110011011111111111001011100111111",
   "110101011010000000101100100100001011111111111101011101110001001011",
   "110101011100000000101100100111100001101011111011000010100000000101",
   "110101011110000000101100101010110111011111111000100111101001101101",
   "110101100000000000101100101110001101011011110110001101001110000100",
   "110101100010000000101100110001100011011111110011110011001101001010",
   "110101100100000000101100110100111001101011110001011001100111000010",
   "110101100110000000101100111000001111111111101111000000011011101100",
   "110101101000000000101100111011100110011011101100100111101011001001",
   "110101101010000000101100111110111100111111101010001111010101011001",
   "110101101100000000101101000010010011101011100111110111011010011111",
   "110101101110000000101101000101101010011111100101011111111010011011",
   "110101110000000000101101001001000001011011100011001000110101001110",
   "110101110010000000101101001100011000011111100000110010001010111001",
   "110101110100000000101101001111101111101011011110011011111011011100",
   "110101110110000000101101010011000110111111011100000110000110111010",
   "110101111000000000101101010110011110011011011001110000101101010011",
   "110101111010000000101101011001110101111111010111011011101110101000",
   "110101111100000000101101011101001101101011010101000111001010111001",
   "110101111110000000101101100000100101011111010010110011000010001001",
   "110110000000000000101101100011111101011011010000011111010100011000",
   "110110000010000000101101100111010101011111001110001100000001100111",
   "110110000100000000101101101010101101101011001011111001001001110111",
   "110110000110000000101101101110000101111111001001100110101101001000",
   "110110001000000000101101110001011110011011000111010100101011011101",
   "110110001010000000101101110100110110111111000101000011000100110110",
   "110110001100000000101101111000001111101011000010110001111001010100",
   "110110001110000000101101111011101000011111000000100001001000110111",
   "110110010000000000101101111111000001011010111110010000110011100010",
   "110110010010000000101110000010011010011110111100000000111001010101",
   "110110010100000000101110000101110011101010111001110001011010010001",
   "110110010110000000101110001001001100111110110111100010010110010111",
   "110110011000000000101110001100100110011010110101010011101101100111",
   "110110011010000000101110001111111111111110110011000101100000000100",
   "110110011100000000101110010011011001101010110000110111101101101110",
   "110110011110000000101110010110110011011110101110101010010110100110",
   "110110100000000000101110011010001101011010101100011101011010101101",
   "110110100010000000101110011101100111011110101010010000111010000011",
   "110110100100000000101110100001000001101010101000000100110100101011",
   "110110100110000000101110100100011011111110100101111001001010100101",
   "110110101000000000101110100111110110011010100011101101111011110010",
   "110110101010000000101110101011010000111110100001100011001000010011",
   "110110101100000000101110101110101011101010011111011000110000001000",
   "110110101110000000101110110010000110011110011101001110110011010100",
   "110110110000000000101110110101100001011010011011000101010001110111",
   "110110110010000000101110111000111100011110011000111100001011110010",
   "110110110100000000101110111100010111101010010110110011100001000110",
   "110110110110000000101110111111110010111110010100101011010001110011",
   "110110111000000000101111000011001110011010010010100011011101111100",
   "110110111010000000101111000110101001111110010000011100000101100001",
   "110110111100000000101111001010000101101010001110010101001000100011",
   "110110111110000000101111001101100001011110001100001110100111000011",
   "110111000000000000101111010000111101011010001010001000100001000001",
   "110111000010000000101111010100011001011110001000000010110110100000",
   "110111000100000000101111010111110101101010000101111101100111100000",
   "110111000110000000101111011011010001111110000011111000110100000010",
   "110111001000000000101111011110101110011010000001110100011100000111",
   "110111001010000000101111100010001010111101111111110000011111110000",
   "110111001100000000101111100101100111101001111101101100111110111101",
   "110111001110000000101111101001000100011101111011101001111001110001",
   "110111010000000000101111101100100001011001111001100111010000001100",
   "110111010010000000101111101111111110011101110111100101000010001111",
   "110111010100000000101111110011011011101001110101100011001111111011",
   "110111010110000000101111110110111000111101110011100001111001010001",
   "110111011000000000101111111010010110011001110001100000111110010001",
   "110111011010000000101111111101110011111101101111100000011110111110",
   "110111011100000000110000000001010001101001101101100000011011011000",
   "110111011110000000110000000100101111011101101011100000110011100000",
   "110111100000000000110000001000001101011001101001100001100111010111",
   "110111100010000000110000001011101011011101100111100010110110111110",
   "110111100100000000110000001111001001101001100101100100100010010110",
   "110111100110000000110000010010100111111101100011100110101001011111",
   "110111101000000000110000010110000110011001100001101001001100011100",
   "110111101010000000110000011001100100111101011111101100001011001101",
   "110111101100000000110000011101000011101001011101101111100101110011",
   "110111101110000000110000100000100010011101011011110011011100001111",
   "110111110000000000110000100100000001011001011001110111101110100010",
   "110111110010000000110000100111100000011101010111111100011100101101",
   "110111110100000000110000101010111111101001010110000001100110110000",
   "110111110110000000110000101110011110111101010100000111001100101110",
   "110111111000000000110000110001111110011001010010001101001110100111",
   "110111111010000000110000110101011101111101010000010011101100011100",
   "110111111100000000110000111000111101101001001110011010100110001110",
   "110111111110000000110000111100011101011101001100100001111011111110",
   "111000000000000000110000111111111101011001001010101001101101101101",
   "111000000010000000110001000011011101011101001000110001111011011100",
   "111000000100000000110001000110111101101001000110111010100101001100",
   "111000000110000000110001001010011101111101000101000011101010111101",
   "111000001000000000110001001101111110011001000011001101001100110010",
   "111000001010000000110001010001011110111101000001010111001010101011",
   "111000001100000000110001010100111111101000111111100001100100101001",
   "111000001110000000110001011000100000011100111101101100011010101101",
   "111000010000000000110001011100000001011000111011110111101100111000",
   "111000010010000000110001011111100010011100111010000011011011001011",
   "111000010100000000110001100011000011101000111000001111100101100111",
   "111000010110000000110001100110100100111100110110011100001100001101",
   "111000011000000000110001101010000110011000110100101001001110111110",
   "111000011010000000110001101101100111111100110010110110101101111010",
   "111000011100000000110001110001001001101000110001000100101001000100",
   "111000011110000000110001110100101011011100101111010011000000011100",
   "111000100000000000110001111000001101011000101101100001110100000011",
   "111000100010000000110001111011101111011100101011110001000011111010",
   "111000100100000000110001111111010001101000101010000000110000000010",
   "111000100110000000110010000010110011111100101000010000111000011100",
   "111000101000000000110010000110010110011000100110100001011101001001",
   "111000101010000000110010001001111000111100100100110010011110001010",
   "111000101100000000110010001101011011101000100011000011111011100000",
   "111000101110000000110010010000111110011100100001010101110101001100",
   "111000110000000000110010010100100001011000011111101000001011001111",
   "111000110010000000110010011000000100011100011101111010111101101010",
   "111000110100000000110010011011100111101000011100001110001100011110",
   "111000110110000000110010011111001010111100011010100001110111101100",
   "111000111000000000110010100010101110011000011000110101111111010101",
   "111000111010000000110010100110010001111100010111001010100011011001",
   "111000111100000000110010101001110101101000010101011111100011111011",
   "111000111110000000110010101101011001011100010011110101000000111011",
   "111001000000000000110010110000111101011000010010001010111010011010",
   "111001000010000000110010110100100001011100010000100001010000011001",
   "111001000100000000110010111000000101101000001110111000000010111001",
   "111001000110000000110010111011101001111100001101001111010001111011",
   "111001001000000000110010111111001110011000001011100110111101100000",
   "111001001010000000110011000010110010111100001001111111000101101001",
   "111001001100000000110011000110010111101000001000010111101010010111",
   "111001001110000000110011001001111100011100000110110000101011101011",
   "111001010000000000110011001101100001011000000101001010001001100110",
   "111001010010000000110011010001000110011100000011100100000100001001",
   "111001010100000000110011010100101011101000000001111110011011010101",
   "111001010110000000110011011000010000111100000000011001001111001011",
   "111001011000000000110011011011110110010111111110110100011111101100",
   "111001011010000000110011011111011011111011111101010000001100111001",
   "111001011100000000110011100011000001100111111011101100010110110011",
   "111001011110000000110011100110100111011011111010001000111101011011",
   "111001100000000000110011101010001101010111111000100110000000110010",
   "111001100010000000110011101101110011011011110111000011100000111001",
   "111001100100000000110011110001011001100111110101100001011101110001",
   "111001100110000000110011110100111111111011110011111111110111011011",
   "111001101000000000110011111000100110010111110010011110101101111000",
   "111001101010000000110011111100001100111011110000111110000001001001",
   "111001101100000000110011111111110011100111101111011101110001001111",
   "111001101110000000110100000011011010011011101101111101111110001100",
   "111001110000000000110100000111000001010111101100011110100111111111",
   "111001110010000000110100001010101000011011101010111111101110101010",
   "111001110100000000110100001110001111100111101001100001010010001110",
   "111001110110000000110100010001110110111011101000000011010010101100",
   "111001111000000000110100010101011110010111100110100101110000000101",
   "111001111010000000110100011001000101111011100101001000101010011010",
   "111001111100000000110100011100101101100111100011101100000001101100",
   "111001111110000000110100100000010101011011100010001111110101111100",
   "111010000000000000110100100011111101010111100000110100000111001011",
   "111010000010000000110100100111100101011011011111011000110101011010",
   "111010000100000000110100101011001101100111011101111110000000101010",
   "111010000110000000110100101110110101111011011100100011101000111100",
   "111010001000000000110100110010011110010111011011001001101110010001",
   "111010001010000000110100110110000110111011011001110000010000101010",
   "111010001100000000110100111001101111100111011000010111010000001001",
   "111010001110000000110100111101011000011011010110111110101100101101",
   "111010010000000000110101000001000001010111010101100110100110011000",
   "111010010010000000110101000100101010011011010100001110111101001011",
   "111010010100000000110101001000010011100111010010110111110001000111",
   "111010010110000000110101001011111100111011010001100001000010001101",
   "111010011000000000110101001111100110010111010000001010110000011110",
   "111010011010000000110101010011001111111011001110110100111011111011",
   "111010011100000000110101010110111001100111001101011111100100100101",
   "111010011110000000110101011010100011011011001100001010101010011110",
   "111010100000000000110101011110001101010111001010110110001101100101",
   "111010100010000000110101100001110111011011001001100010001101111100",
   "111010100100000000110101100101100001100111001000001110101011100100",
   "111010100110000000110101101001001011111011000110111011100110011110",
   "111010101000000000110101101100110110010111000101101000111110101011",
   "111010101010000000110101110000100000111011000100010110110100001100",
   "111010101100000000110101110100001011100111000011000101000111000011",
   "111010101110000000110101110111110110011011000001110011110111001111",
   "111010110000000000110101111011100001010111000000100011000100110010",
   "111010110010000000110101111111001100011010111111010010101111101101",
   "111010110100000000110110000010110111100110111110000010111000000001",
   "111010110110000000110110000110100010111010111100110011011101101111",
   "111010111000000000110110001010001110010110111011100100100000111001",
   "111010111010000000110110001101111001111010111010010110000001011110",
   "111010111100000000110110010001100101100110111001000111111111100000",
   "111010111110000000110110010101010001011010110111111010011011000000",
   "111011000000000000110110011000111101010110110110101101010011111111",
   "111011000010000000110110011100101001011010110101100000101010011111",
   "111011000100000000110110100000010101100110110100010100011110011111",
   "111011000110000000110110100100000001111010110011001000110000000001",
   "111011001000000000110110100111101110010110110001111101011111000110",
   "111011001010000000110110101011011010111010110000110010101011101111",
   "111011001100000000110110101111000111100110101111101000010101111110",
   "111011001110000000110110110010110100011010101110011110011101110010",
   "111011010000000000110110110110100001010110101101010101000011001101",
   "111011010010000000110110111010001110011010101100001100000110010000",
   "111011010100000000110110111101111011100110101011000011100110111101",
   "111011010110000000110111000001101000111010101001111011100101010011",
   "111011011000000000110111000101010110010110101000110100000001010100",
   "111011011010000000110111001001000011111010100111101100111011000001",
   "111011011100000000110111001100110001100110100110100110010010011100",
   "111011011110000000110111010000011111011010100101100000000111100100",
   "111011100000000000110111010100001101010110100100011010011010011011",
   "111011100010000000110111010111111011011010100011010101001011000010",
   "111011100100000000110111011011101001100110100010010000011001011011",
   "111011100110000000110111011111010111111010100001001100000101100101",
   "111011101000000000110111100011000110010110100000001000001111100010",
   "111011101010000000110111100110110100111010011111000100110111010100",
   "111011101100000000110111101010100011100110011110000001111100111010",
   "111011101110000000110111101110010010011010011100111111100000010110",
   "111011110000000000110111110010000001010110011011111101100001101010",
   "111011110010000000110111110101110000011010011010111100000000110101",
   "111011110100000000110111111001011111100110011001111010111101111001",
   "111011110110000000110111111101001110111010011000111010011000111000",
   "111011111000000000111000000000111110010110010111111010010001110001",
   "111011111010000000111000000100101101111010010110111010101000100110",
   "111011111100000000111000001000011101100110010101111011011101011000",
   "111011111110000000111000001100001101011010010100111100110000001001",
   "111100000000000000111000001111111101010110010011111110100000111000",
   "111100000010000000111000010011101101011010010011000000101111101000",
   "111100000100000000111000010111011101100110010010000011011100011000",
   "111100000110000000111000011011001101111010010001000110100111001010",
   "111100001000000000111000011110111110010110010000001010010000000000",
   "111100001010000000111000100010101110111010001111001110010110111001",
   "111100001100000000111000100110011111100110001110010010111011110111",
   "111100001110000000111000101010010000011010001101010111111110111100",
   "111100010000000000111000101110000001010110001100011101100000000111",
   "111100010010000000111000110001110010011010001011100011011111011011",
   "111100010100000000111000110101100011100110001010101001111100110111",
   "111100010110000000111000111001010100111010001001110000111000011101",
   "111100011000000000111000111101000110010110001000111000010010001111",
   "111100011010000000111001000000110111111010001000000000001010001100",
   "111100011100000000111001000100101001100110000111001000100000010111",
   "111100011110000000111001001000011011011010000110010001010100101111",
   "111100100000000000111001001100001101010110000101011010100111010110",
   "111100100010000000111001001111111111011010000100100100011000001110",
   "111100100100000000111001010011110001100110000011101110100111010110",
   "111100100110000000111001010111100011111010000010111001010100110001",
   "111100101000000000111001011011010110010110000010000100100000011110",
   "111100101010000000111001011111001000111010000001010000001010100000",
   "111100101100000000111001100010111011100110000000011100010010110110",
   "111100101110000000111001100110101110011001111111101000111001100011",
   "111100110000000000111001101010100001010101111110110101111110100110",
   "111100110010000000111001101110010100011001111110000011100010000010",
   "111100110100000000111001110010000111100101111101010001100011110110",
   "111100110110000000111001110101111010111001111100100000000100000101",
   "111100111000000000111001111001101110010101111011101111000010101110",
   "111100111010000000111001111101100001111001111010111110011111110100",
   "111100111100000000111010000001010101100101111010001110011011010110",
   "111100111110000000111010000101001001011001111001011110110101010111",
   "111101000000000000111010001000111101010101111000101111101101110110",
   "111101000010000000111010001100110001011001111000000001000100110110",
   "111101000100000000111010010000100101100101110111010010111010010110",
   "111101000110000000111010010100011001111001110110100101001110011001",
   "111101001000000000111010011000001110010101110101111000000000111110",
   "111101001010000000111010011100000010111001110101001011010010001000",
   "111101001100000000111010011111110111100101110100011111000001110110",
   "111101001110000000111010100011101100011001110011110011010000001011",
   "111101010000000000111010100111100001010101110011000111111101000110",
   "111101010010000000111010101011010110011001110010011101001000101010",
   "111101010100000000111010101111001011100101110001110010110010110111",
   "111101010110000000111010110011000000111001110001001000111011101101",
   "111101011000000000111010110110110110010101110000011111100011001111",
   "111101011010000000111010111010101011111001101111110110101001011100",
   "111101011100000000111010111110100001100101101111001110001110010111",
   "111101011110000000111011000010010111011001101110100110010010000000",
   "111101100000000000111011000110001101010101101101111110110100010111",
   "111101100010000000111011001010000011011001101101010111110101011111",
   "111101100100000000111011001101111001100101101100110001010101010111",
   "111101100110000000111011010001101111111001101100001011010100000010",
   "111101101000000000111011010101100110010101101011100101110001100000",
   "111101101010000000111011011001011100111001101011000000101101110001",
   "111101101100000000111011011101010011100101101010011100001000111000",
   "111101101110000000111011100001001010011001101001111000000010110101",
   "111101110000000000111011100101000001010101101001010100011011101000",
   "111101110010000000111011101000111000011001101000110001010011010100",
   "111101110100000000111011101100101111100101101000001110101001111001",
   "111101110110000000111011110000100110111001100111101100011111010111",
   "111101111000000000111011110100011110010101100111001010110011110001",
   "111101111010000000111011111000010101111001100110101001100111000111",
   "111101111100000000111011111100001101100101100110001000111001011001",
   "111101111110000000111100000000000101011001100101101000101010101010",
   "111110000000000000111100000011111101010101100101001000111010111010",
   "111110000010000000111100000111110101011001100100101001101010001001",
   "111110000100000000111100001011101101100101100100001010111000011010",
   "111110000110000000111100001111100101111001100011101100100101101101",
   "111110001000000000111100010011011110010101100011001110110010000011",
   "111110001010000000111100010111010110111001100010110001011101011100",
   "111110001100000000111100011011001111100101100010010100100111111011",
   "111110001110000000111100011111001000011001100001111000010001100000",
   "111110010000000000111100100011000001010101100001011100011010001100",
   "111110010010000000111100100110111010011001100001000001000001111111",
   "111110010100000000111100101010110011100101100000100110001000111100",
   "111110010110000000111100101110101100111001100000001011101111000011",
   "111110011000000000111100110010100110010101011111110001110100010101",
   "111110011010000000111100110110011111111001011111011000011000110011",
   "111110011100000000111100111010011001100101011110111111011100011101",
   "111110011110000000111100111110010011011001011110100110111111010110",
   "111110100000000000111101000010001101010101011110001111000001011110",
   "111110100010000000111101000110000111011001011101110111100010110110",
   "111110100100000000111101001010000001100101011101100000100011011111",
   "111110100110000000111101001101111011111001011101001010000011011001",
   "111110101000000000111101010001110110010101011100110100000010100111",
   "111110101010000000111101010101110000111001011100011110100001001001",
   "111110101100000000111101011001101011100101011100001001011111000000",
   "111110101110000000111101011101100110011001011011110100111100001101",
   "111110110000000000111101100001100001010101011011100000111000110001",
   "111110110010000000111101100101011100011001011011001101010100101101",
   "111110110100000000111101101001010111100101011010111010010000000001",
   "111110110110000000111101101101010010111001011010100111101010110000",
   "111110111000000000111101110001001110010101011010010101100100111010",
   "111110111010000000111101110101001001111001011010000011111110100000",
   "111110111100000000111101111001000101100101011001110010110111100011",
   "111110111110000000111101111101000001011001011001100010010000000100",
   "111111000000000000111110000000111101010101011001010010001000000100",
   "111111000010000000111110000100111001011001011001000010011111100100",
   "111111000100000000111110001000110101100101011000110011010110100101",
   "111111000110000000111110001100110001111001011000100100101101001000",
   "111111001000000000111110010000101110010101011000010110100011001110",
   "111111001010000000111110010100101010111001011000001000111000111000",
   "111111001100000000111110011000100111100101010111111011101110000111",
   "111111001110000000111110011100100100011001010111101111000010111100",
   "111111010000000000111110100000100001010101010111100010110111011000",
   "111111010010000000111110100100011110011001010111010111001011011100",
   "111111010100000000111110101000011011100101010111001011111111001001",
   "111111010110000000111110101100011000111001010111000001010010100000",
   "111111011000000000111110110000010110010101010110110111000101100010",
   "111111011010000000111110110100010011111001010110101101011000010000",
   "111111011100000000111110111000010001100101010110100100001010101011",
   "111111011110000000111110111100001111011001010110011011011100110100",
   "111111100000000000111111000000001101010101010110010011001110101100",
   "111111100010000000111111000100001011011001010110001011100000010100",
   "111111100100000000111111001000001001100101010110000100010001101101",
   "111111100110000000111111001100000111111001010101111101100010111000",
   "111111101000000000111111010000000110010101010101110111010011110110",
   "111111101010000000111111010100000100111001010101110001100100101000",
   "111111101100000000111111011000000011100101010101101100010101001111",
   "111111101110000000111111011100000010011001010101100111100101101100",
   "111111110000000000111111100000000001010101010101100011010110000000",
   "111111110010000000111111100100000000011001010101011111100110001100",
   "111111110100000000111111100111111111100101010101011100010110010010",
   "111111110110000000111111101011111110111001010101011001100110010001",
   "111111111000000000111111101111111110010101010101010111010110001011",
   "111111111010000000111111110011111101111001010101010101100110000001",
   "111111111100000000111111110111111101100101010101010100010101110100",
   "111111111110000000111111111011111101011001010101010011100101100101",
      others => (others => '0'));
      	begin 
      return tmp;
      end init_rom;
	signal rom : memory_t := init_rom;
   signal Y0 :  std_logic_vector(65 downto 0);
begin
	process(clk)
   begin
   if(rising_edge(clk)) then
   	Y0 <= rom(  TO_INTEGER(unsigned(X))  );
   end if;
   end process;
    Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_83_f400_uid137
--                     (IntAdderClassical_83_f400_uid139)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_83_f400_uid137 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(82 downto 0);
          Y : in  std_logic_vector(82 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(82 downto 0)   );
end entity;

architecture arch of IntAdder_83_f400_uid137 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_83_f400_uid144
--                     (IntAdderClassical_83_f400_uid146)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_83_f400_uid144 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(82 downto 0);
          Y : in  std_logic_vector(82 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(82 downto 0)   );
end entity;

architecture arch of IntAdder_83_f400_uid144 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                   KCMTable_6_49946518145322874_unsigned
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity KCMTable_6_49946518145322874_unsigned is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(61 downto 0)   );
end entity;

architecture arch of KCMTable_6_49946518145322874_unsigned is
begin
  with X select  Y <= 
   "00000000000000000000000000000000000000000000000000000000000000" when "000000",
   "00000010110001011100100001011111110111110100011100111101111010" when "000001",
   "00000101100010111001000010111111101111101000111001111011110100" when "000010",
   "00001000010100010101100100011111100111011101010110111001101110" when "000011",
   "00001011000101110010000101111111011111010001110011110111101000" when "000100",
   "00001101110111001110100111011111010111000110010000110101100010" when "000101",
   "00010000101000101011001000111111001110111010101101110011011100" when "000110",
   "00010011011010000111101010011111000110101111001010110001010110" when "000111",
   "00010110001011100100001011111110111110100011100111101111010000" when "001000",
   "00011000111101000000101101011110110110011000000100101101001010" when "001001",
   "00011011101110011101001110111110101110001100100001101011000100" when "001010",
   "00011110011111111001110000011110100110000000111110101000111110" when "001011",
   "00100001010001010110010001111110011101110101011011100110111000" when "001100",
   "00100100000010110010110011011110010101101001111000100100110010" when "001101",
   "00100110110100001111010100111110001101011110010101100010101100" when "001110",
   "00101001100101101011110110011110000101010010110010100000100110" when "001111",
   "00101100010111001000010111111101111101000111001111011110100000" when "010000",
   "00101111001000100100111001011101110100111011101100011100011010" when "010001",
   "00110001111010000001011010111101101100110000001001011010010100" when "010010",
   "00110100101011011101111100011101100100100100100110011000001110" when "010011",
   "00110111011100111010011101111101011100011001000011010110001000" when "010100",
   "00111010001110010110111111011101010100001101100000010100000010" when "010101",
   "00111100111111110011100000111101001100000001111101010001111100" when "010110",
   "00111111110001010000000010011101000011110110011010001111110110" when "010111",
   "01000010100010101100100011111100111011101010110111001101110000" when "011000",
   "01000101010100001001000101011100110011011111010100001011101010" when "011001",
   "01001000000101100101100110111100101011010011110001001001100100" when "011010",
   "01001010110111000010001000011100100011001000001110000111011110" when "011011",
   "01001101101000011110101001111100011010111100101011000101011000" when "011100",
   "01010000011001111011001011011100010010110001001000000011010010" when "011101",
   "01010011001011010111101100111100001010100101100101000001001100" when "011110",
   "01010101111100110100001110011100000010011010000001111111000110" when "011111",
   "01011000101110010000101111111011111010001110011110111101000000" when "100000",
   "01011011011111101101010001011011110010000010111011111010111010" when "100001",
   "01011110010001001001110010111011101001110111011000111000110100" when "100010",
   "01100001000010100110010100011011100001101011110101110110101110" when "100011",
   "01100011110100000010110101111011011001100000010010110100101000" when "100100",
   "01100110100101011111010111011011010001010100101111110010100010" when "100101",
   "01101001010110111011111000111011001001001001001100110000011100" when "100110",
   "01101100001000011000011010011011000000111101101001101110010110" when "100111",
   "01101110111001110100111011111010111000110010000110101100010000" when "101000",
   "01110001101011010001011101011010110000100110100011101010001010" when "101001",
   "01110100011100101101111110111010101000011011000000101000000100" when "101010",
   "01110111001110001010100000011010100000001111011101100101111110" when "101011",
   "01111001111111100111000001111010011000000011111010100011111000" when "101100",
   "01111100110001000011100011011010001111111000010111100001110010" when "101101",
   "01111111100010100000000100111010000111101100110100011111101100" when "101110",
   "10000010010011111100100110011001111111100001010001011101100110" when "101111",
   "10000101000101011001000111111001110111010101101110011011100000" when "110000",
   "10000111110110110101101001011001101111001010001011011001011010" when "110001",
   "10001010101000010010001010111001100110111110101000010111010100" when "110010",
   "10001101011001101110101100011001011110110011000101010101001110" when "110011",
   "10010000001011001011001101111001010110100111100010010011001000" when "110100",
   "10010010111100100111101111011001001110011011111111010001000010" when "110101",
   "10010101101110000100010000111001000110010000011100001110111100" when "110110",
   "10011000011111100000110010011000111110000100111001001100110110" when "110111",
   "10011011010000111101010011111000110101111001010110001010110000" when "111000",
   "10011110000010011001110101011000101101101101110011001000101010" when "111001",
   "10100000110011110110010110111000100101100010010000000110100100" when "111010",
   "10100011100101010010111000011000011101010110101101000100011110" when "111011",
   "10100110010110101111011001111000010101001011001010000010011000" when "111100",
   "10101001001000001011111011011000001100111111100111000000010010" when "111101",
   "10101011111001101000011100111000000100110100000011111110001100" when "111110",
   "10101110101011000100111110010111111100101000100000111100000110" when "111111",
   "--------------------------------------------------------------" when others;
end architecture;

--------------------------------------------------------------------------------
--                   KCMTable_5_49946518145322874_unsigned
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity KCMTable_5_49946518145322874_unsigned is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(60 downto 0)   );
end entity;

architecture arch of KCMTable_5_49946518145322874_unsigned is
begin
  with X select  Y <= 
   "0000000000000000000000000000000000000000000000000000000000000" when "00000",
   "0000010110001011100100001011111110111110100011100111101111010" when "00001",
   "0000101100010111001000010111111101111101000111001111011110100" when "00010",
   "0001000010100010101100100011111100111011101010110111001101110" when "00011",
   "0001011000101110010000101111111011111010001110011110111101000" when "00100",
   "0001101110111001110100111011111010111000110010000110101100010" when "00101",
   "0010000101000101011001000111111001110111010101101110011011100" when "00110",
   "0010011011010000111101010011111000110101111001010110001010110" when "00111",
   "0010110001011100100001011111110111110100011100111101111010000" when "01000",
   "0011000111101000000101101011110110110011000000100101101001010" when "01001",
   "0011011101110011101001110111110101110001100100001101011000100" when "01010",
   "0011110011111111001110000011110100110000000111110101000111110" when "01011",
   "0100001010001010110010001111110011101110101011011100110111000" when "01100",
   "0100100000010110010110011011110010101101001111000100100110010" when "01101",
   "0100110110100001111010100111110001101011110010101100010101100" when "01110",
   "0101001100101101011110110011110000101010010110010100000100110" when "01111",
   "0101100010111001000010111111101111101000111001111011110100000" when "10000",
   "0101111001000100100111001011101110100111011101100011100011010" when "10001",
   "0110001111010000001011010111101101100110000001001011010010100" when "10010",
   "0110100101011011101111100011101100100100100100110011000001110" when "10011",
   "0110111011100111010011101111101011100011001000011010110001000" when "10100",
   "0111010001110010110111111011101010100001101100000010100000010" when "10101",
   "0111100111111110011100000111101001100000001111101010001111100" when "10110",
   "0111111110001010000000010011101000011110110011010001111110110" when "10111",
   "1000010100010101100100011111100111011101010110111001101110000" when "11000",
   "1000101010100001001000101011100110011011111010100001011101010" when "11001",
   "1001000000101100101100110111100101011010011110001001001100100" when "11010",
   "1001010110111000010001000011100100011001000001110000111011110" when "11011",
   "1001101101000011110101001111100011010111100101011000101011000" when "11100",
   "1010000011001111011001011011100010010110001001000000011010010" when "11101",
   "1010011001011010111101100111100001010100101100101000001001100" when "11110",
   "1010101111100110100001110011100000010011010000001111111000110" when "11111",
   "-------------------------------------------------------------" when others;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_61_f400_uid156
--                     (IntAdderClassical_61_f400_uid158)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_61_f400_uid156 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(60 downto 0);
          Y : in  std_logic_vector(60 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(60 downto 0)   );
end entity;

architecture arch of IntAdder_61_f400_uid156 is
signal X_d1 :  std_logic_vector(60 downto 0);
signal Y_d1 :  std_logic_vector(60 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
    R <= X_d1 + Y_d1 + Cin_d1;
end architecture;

--------------------------------------------------------------------------------
--                  IntIntKCM_11_49946518145322874_unsigned
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2009,2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntIntKCM_11_49946518145322874_unsigned is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          R : out  std_logic_vector(66 downto 0)   );
end entity;

architecture arch of IntIntKCM_11_49946518145322874_unsigned is
   component IntAdder_61_f400_uid156 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(60 downto 0);
             Y : in  std_logic_vector(60 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(60 downto 0)   );
   end component;

   component KCMTable_5_49946518145322874_unsigned is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(60 downto 0)   );
   end component;

   component KCMTable_6_49946518145322874_unsigned is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(61 downto 0)   );
   end component;

signal d0 :  std_logic_vector(5 downto 0);
signal pp0, pp0_d1 :  std_logic_vector(61 downto 0);
signal d1 :  std_logic_vector(4 downto 0);
signal pp1 :  std_logic_vector(60 downto 0);
signal addOp0 :  std_logic_vector(60 downto 0);
signal addOp1 :  std_logic_vector(60 downto 0);
signal OutRes :  std_logic_vector(60 downto 0);
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of KCMTable_5_49946518145322874_unsigned: component is "yes";
attribute rom_extract of KCMTable_6_49946518145322874_unsigned: component is "yes";
attribute rom_style of KCMTable_5_49946518145322874_unsigned: component is "distributed";
attribute rom_style of KCMTable_6_49946518145322874_unsigned: component is "distributed";
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            pp0_d1 <=  pp0;
         end if;
      end process;
   d0 <= X(5 downto 0);
   KCMTable_0: KCMTable_6_49946518145322874_unsigned  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => d0,
                 Y => pp0);
   d1 <= X(10 downto 6);
   KCMTable_1: KCMTable_5_49946518145322874_unsigned  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => d1,
                 Y => pp1);
   addOp0 <= (60 downto 56 => '0') & pp0(61 downto 6) & "";
   addOp1 <= pp1(60 downto 0) & "";
   Result_Adder: IntAdder_61_f400_uid156  -- pipelineDepth=1 maxInDelay=1.6493e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => '0',
                 R => OutRes,
                 X => addOp0,
                 Y => addOp1);
   ----------------Synchro barrier, entering cycle 1----------------
   R <= OutRes & pp0_d1(5 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_94_f400_uid164
--                     (IntAdderClassical_94_f400_uid166)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_94_f400_uid164 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(93 downto 0);
          Y : in  std_logic_vector(93 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(93 downto 0)   );
end entity;

architecture arch of IntAdder_94_f400_uid164 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                  LZCShifter_94_to_83_counting_128_uid171
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_94_to_83_counting_128_uid171 is
   port ( clk, rst : in std_logic;
          I : in  std_logic_vector(93 downto 0);
          Count : out  std_logic_vector(6 downto 0);
          O : out  std_logic_vector(82 downto 0)   );
end entity;

architecture arch of LZCShifter_94_to_83_counting_128_uid171 is
signal level7, level7_d1 :  std_logic_vector(93 downto 0);
signal count6, count6_d1, count6_d2, count6_d3 : std_logic;
signal level6 :  std_logic_vector(93 downto 0);
signal count5, count5_d1, count5_d2, count5_d3 : std_logic;
signal level5, level5_d1 :  std_logic_vector(93 downto 0);
signal count4, count4_d1, count4_d2 : std_logic;
signal level4 :  std_logic_vector(93 downto 0);
signal count3, count3_d1, count3_d2 : std_logic;
signal level3, level3_d1 :  std_logic_vector(89 downto 0);
signal count2, count2_d1 : std_logic;
signal level2 :  std_logic_vector(85 downto 0);
signal count1, count1_d1 : std_logic;
signal level1, level1_d1 :  std_logic_vector(83 downto 0);
signal count0 : std_logic;
signal level0 :  std_logic_vector(82 downto 0);
signal sCount :  std_logic_vector(6 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            level7_d1 <=  level7;
            count6_d1 <=  count6;
            count6_d2 <=  count6_d1;
            count6_d3 <=  count6_d2;
            count5_d1 <=  count5;
            count5_d2 <=  count5_d1;
            count5_d3 <=  count5_d2;
            level5_d1 <=  level5;
            count4_d1 <=  count4;
            count4_d2 <=  count4_d1;
            count3_d1 <=  count3;
            count3_d2 <=  count3_d1;
            level3_d1 <=  level3;
            count2_d1 <=  count2;
            count1_d1 <=  count1;
            level1_d1 <=  level1;
         end if;
      end process;
   level7 <= I ;
   ----------------Synchro barrier, entering cycle 1----------------
   count6<= '1' when level7_d1(93 downto 30) = (93 downto 30=>'0') else '0';
   level6<= level7_d1(93 downto 0) when count6='0' else level7_d1(29 downto 0) & (63 downto 0 => '0');

   count5<= '1' when level6(93 downto 62) = (93 downto 62=>'0') else '0';
   level5<= level6(93 downto 0) when count5='0' else level6(61 downto 0) & (31 downto 0 => '0');

   ----------------Synchro barrier, entering cycle 2----------------
   count4<= '1' when level5_d1(93 downto 78) = (93 downto 78=>'0') else '0';
   level4<= level5_d1(93 downto 0) when count4='0' else level5_d1(77 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(93 downto 86) = (93 downto 86=>'0') else '0';
   level3<= level4(93 downto 4) when count3='0' else level4(85 downto 0) & (3 downto 0 => '0');

   ----------------Synchro barrier, entering cycle 3----------------
   count2<= '1' when level3_d1(89 downto 86) = (89 downto 86=>'0') else '0';
   level2<= level3_d1(89 downto 4) when count2='0' else level3_d1(85 downto 0);

   count1<= '1' when level2(85 downto 84) = (85 downto 84=>'0') else '0';
   level1<= level2(85 downto 2) when count1='0' else level2(83 downto 0);

   ----------------Synchro barrier, entering cycle 4----------------
   count0<= '1' when level1_d1(83 downto 83) = (83 downto 83=>'0') else '0';
   level0<= level1_d1(83 downto 1) when count0='0' else level1_d1(82 downto 0);

   O <= level0;
   sCount <= count6_d3 & count5_d3 & count4_d2 & count3_d2 & count2_d1 & count1_d1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                      RightShifter_31_by_max_30_uid174
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifter_31_by_max_30_uid174 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(30 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(60 downto 0)   );
end entity;

architecture arch of RightShifter_31_by_max_30_uid174 is
signal level0, level0_d1 :  std_logic_vector(30 downto 0);
signal ps, ps_d1 :  std_logic_vector(4 downto 0);
signal level1 :  std_logic_vector(31 downto 0);
signal level2 :  std_logic_vector(33 downto 0);
signal level3 :  std_logic_vector(37 downto 0);
signal level4 :  std_logic_vector(45 downto 0);
signal level5 :  std_logic_vector(61 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            level0_d1 <=  level0;
            ps_d1 <=  ps;
         end if;
      end process;
   level0<= X;
   ps<= S;
   ----------------Synchro barrier, entering cycle 1----------------
   level1<=  (0 downto 0 => '0') & level0_d1 when ps_d1(0) = '1' else    level0_d1 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps_d1(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps_d1(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps_d1(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps_d1(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(61 downto 1);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_58_f400_uid177
--                     (IntAdderClassical_58_f400_uid179)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_58_f400_uid177 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(57 downto 0);
          Y : in  std_logic_vector(57 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(57 downto 0)   );
end entity;

architecture arch of IntAdder_58_f400_uid177 is
signal X_d1 :  std_logic_vector(57 downto 0);
signal Y_d1 :  std_logic_vector(57 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
    R <= X_d1 + Y_d1 + Cin_d1;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_63_f400_uid184
--                    (IntAdderAlternative_63_f400_uid188)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_63_f400_uid184 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(62 downto 0);
          Y : in  std_logic_vector(62 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(62 downto 0)   );
end entity;

architecture arch of IntAdder_63_f400_uid184 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                                   LPR_Ln
--                            (FPLog_11_52_0_400)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, C. Klein  (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LPR_Ln is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of LPR_Ln is
   component IntAdder_56_f400_uid105 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(55 downto 0);
             Y : in  std_logic_vector(55 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(55 downto 0)   );
   end component;

   component IntAdder_56_f400_uid88 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(55 downto 0);
             Y : in  std_logic_vector(55 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(55 downto 0)   );
   end component;

   component IntAdder_56_f400_uid95 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(55 downto 0);
             Y : in  std_logic_vector(55 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(55 downto 0)   );
   end component;

   component IntAdder_58_f400_uid177 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(57 downto 0);
             Y : in  std_logic_vector(57 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(57 downto 0)   );
   end component;

   component IntAdder_63_f400_uid184 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(62 downto 0);
             Y : in  std_logic_vector(62 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(62 downto 0)   );
   end component;

   component IntAdder_66_f400_uid53 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(65 downto 0);
             Y : in  std_logic_vector(65 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(65 downto 0)   );
   end component;

   component IntAdder_66_f400_uid60 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(65 downto 0);
             Y : in  std_logic_vector(65 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(65 downto 0)   );
   end component;

   component IntAdder_83_f400_uid128 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(82 downto 0);
             Y : in  std_logic_vector(82 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(82 downto 0)   );
   end component;

   component IntAdder_83_f400_uid137 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(82 downto 0);
             Y : in  std_logic_vector(82 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(82 downto 0)   );
   end component;

   component IntAdder_83_f400_uid144 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(82 downto 0);
             Y : in  std_logic_vector(82 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(82 downto 0)   );
   end component;

   component IntAdder_94_f400_uid164 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(93 downto 0);
             Y : in  std_logic_vector(93 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(93 downto 0)   );
   end component;

   component IntIntKCM_11_49946518145322874_unsigned is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             R : out  std_logic_vector(66 downto 0)   );
   end component;

   component IntMultiplier_UsingDSP_11_49_0_unsigned_uid67 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             Y : in  std_logic_vector(48 downto 0);
             R : out  std_logic_vector(59 downto 0)   );
   end component;

   component IntMultiplier_UsingDSP_12_54_0_unsigned_uid11 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(11 downto 0);
             Y : in  std_logic_vector(53 downto 0);
             R : out  std_logic_vector(65 downto 0)   );
   end component;

   component IntMultiplier_UsingDSP_9_55_0_unsigned_uid32 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(8 downto 0);
             Y : in  std_logic_vector(54 downto 0);
             R : out  std_logic_vector(63 downto 0)   );
   end component;

   component IntSquarer_31_uid102 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(30 downto 0);
             R : out  std_logic_vector(61 downto 0)   );
   end component;

   component InvTable_0_11_12 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             Y : out  std_logic_vector(11 downto 0)   );
   end component;

   component LZCShifter_94_to_83_counting_128_uid171 is
      port ( clk, rst : in std_logic;
             I : in  std_logic_vector(93 downto 0);
             Count : out  std_logic_vector(6 downto 0);
             O : out  std_logic_vector(82 downto 0)   );
   end component;

   component LZOC_52_6_uid3 is
      port ( clk, rst : in std_logic;
             I : in  std_logic_vector(51 downto 0);
             OZB : in std_logic;
             O : out  std_logic_vector(5 downto 0)   );
   end component;

   component LeftShifter_27_by_max_27_uid6 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(26 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(53 downto 0)   );
   end component;

   component LogTable_0_11_83 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             Y : out  std_logic_vector(82 downto 0)   );
   end component;

   component LogTable_1_9_74 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(73 downto 0)   );
   end component;

   component LogTable_2_11_66 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             Y : out  std_logic_vector(65 downto 0)   );
   end component;

   component RightShifter_31_by_max_30_uid174 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(30 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(60 downto 0)   );
   end component;

signal XExnSgn, XExnSgn_d1, XExnSgn_d2, XExnSgn_d3, XExnSgn_d4, XExnSgn_d5, XExnSgn_d6, XExnSgn_d7, XExnSgn_d8, XExnSgn_d9, XExnSgn_d10, XExnSgn_d11, XExnSgn_d12, XExnSgn_d13, XExnSgn_d14, XExnSgn_d15, XExnSgn_d16, XExnSgn_d17 :  std_logic_vector(2 downto 0);
signal FirstBit : std_logic;
signal Y0, Y0_d1, Y0_d2 :  std_logic_vector(53 downto 0);
signal Y0h :  std_logic_vector(51 downto 0);
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11, sR_d12, sR_d13, sR_d14, sR_d15, sR_d16, sR_d17 : std_logic;
signal absZ0, absZ0_d1, absZ0_d2, absZ0_d3 :  std_logic_vector(26 downto 0);
signal E :  std_logic_vector(10 downto 0);
signal absE, absE_d1, absE_d2, absE_d3, absE_d4, absE_d5, absE_d6, absE_d7, absE_d8, absE_d9, absE_d10 :  std_logic_vector(10 downto 0);
signal EeqZero, EeqZero_d1, EeqZero_d2, EeqZero_d3 : std_logic;
signal lzo, lzo_d1, lzo_d2, lzo_d3, lzo_d4, lzo_d5, lzo_d6, lzo_d7, lzo_d8, lzo_d9, lzo_d10, lzo_d11, lzo_d12 :  std_logic_vector(5 downto 0);
signal pfinal_s :  std_logic_vector(5 downto 0);
signal shiftval :  std_logic_vector(6 downto 0);
signal shiftvalinL :  std_logic_vector(4 downto 0);
signal shiftvalinR, shiftvalinR_d1, shiftvalinR_d2, shiftvalinR_d3, shiftvalinR_d4, shiftvalinR_d5, shiftvalinR_d6, shiftvalinR_d7, shiftvalinR_d8, shiftvalinR_d9 :  std_logic_vector(4 downto 0);
signal doRR, doRR_d1, doRR_d2, doRR_d3 : std_logic;
signal small, small_d1, small_d2, small_d3, small_d4, small_d5, small_d6, small_d7, small_d8, small_d9, small_d10, small_d11, small_d12, small_d13, small_d14 : std_logic;
signal small_absZ0_normd_full :  std_logic_vector(53 downto 0);
signal small_absZ0_normd, small_absZ0_normd_d1, small_absZ0_normd_d2, small_absZ0_normd_d3, small_absZ0_normd_d4, small_absZ0_normd_d5, small_absZ0_normd_d6, small_absZ0_normd_d7, small_absZ0_normd_d8, small_absZ0_normd_d9 :  std_logic_vector(26 downto 0);
signal A0, A0_d1, A0_d2, A0_d3, A0_d4, A0_d5, A0_d6, A0_d7 :  std_logic_vector(10 downto 0);
signal InvA0 :  std_logic_vector(11 downto 0);
signal P0 :  std_logic_vector(65 downto 0);
signal Z1 :  std_logic_vector(54 downto 0);
signal A1, A1_d1, A1_d2, A1_d3, A1_d4 :  std_logic_vector(8 downto 0);
signal B1 :  std_logic_vector(45 downto 0);
signal ZM1 :  std_logic_vector(54 downto 0);
signal P1 :  std_logic_vector(63 downto 0);
signal Y1 :  std_logic_vector(64 downto 0);
signal EiY1 :  std_logic_vector(65 downto 0);
signal addXIter1 :  std_logic_vector(65 downto 0);
signal EiYPB1, EiYPB1_d1 :  std_logic_vector(65 downto 0);
signal Pp1 :  std_logic_vector(65 downto 0);
signal Z2 :  std_logic_vector(65 downto 0);
signal A2, A2_d1, A2_d2, A2_d3, A2_d4, A2_d5 :  std_logic_vector(10 downto 0);
signal B2 :  std_logic_vector(54 downto 0);
signal ZM2 :  std_logic_vector(48 downto 0);
signal P2 :  std_logic_vector(59 downto 0);
signal Y2 :  std_logic_vector(83 downto 0);
signal EiY2 :  std_logic_vector(55 downto 0);
signal addXIter2 :  std_logic_vector(55 downto 0);
signal EiYPB2 :  std_logic_vector(55 downto 0);
signal Pp2 :  std_logic_vector(55 downto 0);
signal Z3 :  std_logic_vector(55 downto 0);
signal Zfinal, Zfinal_d1, Zfinal_d2, Zfinal_d3, Zfinal_d4 :  std_logic_vector(55 downto 0);
signal squarerIn :  std_logic_vector(30 downto 0);
signal Z2o2_full :  std_logic_vector(61 downto 0);
signal Z2o2_full_dummy, Z2o2_full_dummy_d1, Z2o2_full_dummy_d2 :  std_logic_vector(61 downto 0);
signal Z2o2_normal :  std_logic_vector(27 downto 0);
signal addFinalLog1pY :  std_logic_vector(55 downto 0);
signal Log1p_normal, Log1p_normal_d1 :  std_logic_vector(55 downto 0);
signal L0 :  std_logic_vector(82 downto 0);
signal S1 :  std_logic_vector(82 downto 0);
signal L1 :  std_logic_vector(73 downto 0);
signal sopX1 :  std_logic_vector(82 downto 0);
signal S2, S2_d1, S2_d2 :  std_logic_vector(82 downto 0);
signal L2 :  std_logic_vector(65 downto 0);
signal sopX2 :  std_logic_vector(82 downto 0);
signal S3, S3_d1 :  std_logic_vector(82 downto 0);
signal almostLog :  std_logic_vector(82 downto 0);
signal adderLogF_normalY :  std_logic_vector(82 downto 0);
signal LogF_normal :  std_logic_vector(82 downto 0);
signal absELog2 :  std_logic_vector(66 downto 0);
signal absELog2_pad :  std_logic_vector(93 downto 0);
signal LogF_normal_pad, LogF_normal_pad_d1 :  std_logic_vector(93 downto 0);
signal lnaddX, lnaddX_d1 :  std_logic_vector(93 downto 0);
signal lnaddY :  std_logic_vector(93 downto 0);
signal Log_normal :  std_logic_vector(93 downto 0);
signal E_normal :  std_logic_vector(6 downto 0);
signal Log_normal_normd, Log_normal_normd_d1 :  std_logic_vector(82 downto 0);
signal Z2o2_small_bs :  std_logic_vector(30 downto 0);
signal Z2o2_small_s :  std_logic_vector(60 downto 0);
signal Z2o2_small :  std_logic_vector(57 downto 0);
signal Z_small :  std_logic_vector(57 downto 0);
signal Log_smallY :  std_logic_vector(57 downto 0);
signal nsRCin : std_logic;
signal Log_small, Log_small_d1 :  std_logic_vector(57 downto 0);
signal E0_sub, E0_sub_d1 :  std_logic_vector(1 downto 0);
signal ufl, ufl_d1, ufl_d2, ufl_d3 : std_logic;
signal E_small, E_small_d1 :  std_logic_vector(10 downto 0);
signal Log_small_normd, Log_small_normd_d1, Log_small_normd_d2 :  std_logic_vector(55 downto 0);
signal E0offset :  std_logic_vector(10 downto 0);
signal ER :  std_logic_vector(10 downto 0);
signal Log_g :  std_logic_vector(55 downto 0);
signal round : std_logic;
signal fraX :  std_logic_vector(62 downto 0);
signal fraY :  std_logic_vector(62 downto 0);
signal EFR, EFR_d1 :  std_logic_vector(62 downto 0);
constant g: positive := 4;
constant log2wF: positive := 6;
constant pfinal: positive := 27;
constant sfinal: positive := 56;
constant targetprec: positive := 83;
constant wE: positive := 11;
constant wF: positive := 52;
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of InvTable_0_11_12: component is "yes";
attribute rom_style of InvTable_0_11_12: component is "block";
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            XExnSgn_d1 <=  XExnSgn;
            XExnSgn_d2 <=  XExnSgn_d1;
            XExnSgn_d3 <=  XExnSgn_d2;
            XExnSgn_d4 <=  XExnSgn_d3;
            XExnSgn_d5 <=  XExnSgn_d4;
            XExnSgn_d6 <=  XExnSgn_d5;
            XExnSgn_d7 <=  XExnSgn_d6;
            XExnSgn_d8 <=  XExnSgn_d7;
            XExnSgn_d9 <=  XExnSgn_d8;
            XExnSgn_d10 <=  XExnSgn_d9;
            XExnSgn_d11 <=  XExnSgn_d10;
            XExnSgn_d12 <=  XExnSgn_d11;
            XExnSgn_d13 <=  XExnSgn_d12;
            XExnSgn_d14 <=  XExnSgn_d13;
            XExnSgn_d15 <=  XExnSgn_d14;
            XExnSgn_d16 <=  XExnSgn_d15;
            XExnSgn_d17 <=  XExnSgn_d16;
            Y0_d1 <=  Y0;
            Y0_d2 <=  Y0_d1;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            sR_d12 <=  sR_d11;
            sR_d13 <=  sR_d12;
            sR_d14 <=  sR_d13;
            sR_d15 <=  sR_d14;
            sR_d16 <=  sR_d15;
            sR_d17 <=  sR_d16;
            absZ0_d1 <=  absZ0;
            absZ0_d2 <=  absZ0_d1;
            absZ0_d3 <=  absZ0_d2;
            absE_d1 <=  absE;
            absE_d2 <=  absE_d1;
            absE_d3 <=  absE_d2;
            absE_d4 <=  absE_d3;
            absE_d5 <=  absE_d4;
            absE_d6 <=  absE_d5;
            absE_d7 <=  absE_d6;
            absE_d8 <=  absE_d7;
            absE_d9 <=  absE_d8;
            absE_d10 <=  absE_d9;
            EeqZero_d1 <=  EeqZero;
            EeqZero_d2 <=  EeqZero_d1;
            EeqZero_d3 <=  EeqZero_d2;
            lzo_d1 <=  lzo;
            lzo_d2 <=  lzo_d1;
            lzo_d3 <=  lzo_d2;
            lzo_d4 <=  lzo_d3;
            lzo_d5 <=  lzo_d4;
            lzo_d6 <=  lzo_d5;
            lzo_d7 <=  lzo_d6;
            lzo_d8 <=  lzo_d7;
            lzo_d9 <=  lzo_d8;
            lzo_d10 <=  lzo_d9;
            lzo_d11 <=  lzo_d10;
            lzo_d12 <=  lzo_d11;
            shiftvalinR_d1 <=  shiftvalinR;
            shiftvalinR_d2 <=  shiftvalinR_d1;
            shiftvalinR_d3 <=  shiftvalinR_d2;
            shiftvalinR_d4 <=  shiftvalinR_d3;
            shiftvalinR_d5 <=  shiftvalinR_d4;
            shiftvalinR_d6 <=  shiftvalinR_d5;
            shiftvalinR_d7 <=  shiftvalinR_d6;
            shiftvalinR_d8 <=  shiftvalinR_d7;
            shiftvalinR_d9 <=  shiftvalinR_d8;
            doRR_d1 <=  doRR;
            doRR_d2 <=  doRR_d1;
            doRR_d3 <=  doRR_d2;
            small_d1 <=  small;
            small_d2 <=  small_d1;
            small_d3 <=  small_d2;
            small_d4 <=  small_d3;
            small_d5 <=  small_d4;
            small_d6 <=  small_d5;
            small_d7 <=  small_d6;
            small_d8 <=  small_d7;
            small_d9 <=  small_d8;
            small_d10 <=  small_d9;
            small_d11 <=  small_d10;
            small_d12 <=  small_d11;
            small_d13 <=  small_d12;
            small_d14 <=  small_d13;
            small_absZ0_normd_d1 <=  small_absZ0_normd;
            small_absZ0_normd_d2 <=  small_absZ0_normd_d1;
            small_absZ0_normd_d3 <=  small_absZ0_normd_d2;
            small_absZ0_normd_d4 <=  small_absZ0_normd_d3;
            small_absZ0_normd_d5 <=  small_absZ0_normd_d4;
            small_absZ0_normd_d6 <=  small_absZ0_normd_d5;
            small_absZ0_normd_d7 <=  small_absZ0_normd_d6;
            small_absZ0_normd_d8 <=  small_absZ0_normd_d7;
            small_absZ0_normd_d9 <=  small_absZ0_normd_d8;
            A0_d1 <=  A0;
            A0_d2 <=  A0_d1;
            A0_d3 <=  A0_d2;
            A0_d4 <=  A0_d3;
            A0_d5 <=  A0_d4;
            A0_d6 <=  A0_d5;
            A0_d7 <=  A0_d6;
            A1_d1 <=  A1;
            A1_d2 <=  A1_d1;
            A1_d3 <=  A1_d2;
            A1_d4 <=  A1_d3;
            EiYPB1_d1 <=  EiYPB1;
            A2_d1 <=  A2;
            A2_d2 <=  A2_d1;
            A2_d3 <=  A2_d2;
            A2_d4 <=  A2_d3;
            A2_d5 <=  A2_d4;
            Zfinal_d1 <=  Zfinal;
            Zfinal_d2 <=  Zfinal_d1;
            Zfinal_d3 <=  Zfinal_d2;
            Zfinal_d4 <=  Zfinal_d3;
            Z2o2_full_dummy_d1 <=  Z2o2_full_dummy;
            Z2o2_full_dummy_d2 <=  Z2o2_full_dummy_d1;
            Log1p_normal_d1 <=  Log1p_normal;
            S2_d1 <=  S2;
            S2_d2 <=  S2_d1;
            S3_d1 <=  S3;
            LogF_normal_pad_d1 <=  LogF_normal_pad;
            lnaddX_d1 <=  lnaddX;
            Log_normal_normd_d1 <=  Log_normal_normd;
            Log_small_d1 <=  Log_small;
            E0_sub_d1 <=  E0_sub;
            ufl_d1 <=  ufl;
            ufl_d2 <=  ufl_d1;
            ufl_d3 <=  ufl_d2;
            E_small_d1 <=  E_small;
            Log_small_normd_d1 <=  Log_small_normd;
            Log_small_normd_d2 <=  Log_small_normd_d1;
            EFR_d1 <=  EFR;
         end if;
      end process;
   XExnSgn <=  X(wE+wF+2 downto wE+wF);
   FirstBit <=  X(wF-1);
   Y0 <= "1" & X(wF-1 downto 0) & "0" when FirstBit = '0' else "01" & X(wF-1 downto 0);
   Y0h <= Y0(wF downto 1);
   -- Sign of the result;
   sR <= '0'   when  (X(wE+wF-1 downto wF) = ('0' & (wE-2 downto 0 => '1')))  -- binade [1..2)
     else not X(wE+wF-1);                -- MSB of exponent
   absZ0 <=   Y0(wF-pfinal+1 downto 0)          when (sR='0') else
             ((wF-pfinal+1 downto 0 => '0') - Y0(wF-pfinal+1 downto 0));
   E <= (X(wE+wF-1 downto wF)) - ("0" & (wE-2 downto 1 => '1') & (not FirstBit));
   absE <= ((wE-1 downto 0 => '0') - E)   when sR = '1' else E;
   EeqZero <= '1' when E=(wE-1 downto 0 => '0') else '0';
   ---------------- cycle 0----------------
   lzoc1: LZOC_52_6_uid3  -- pipelineDepth=3 maxInDelay=3.85e-10
      port map ( clk  => clk,
                 rst  => rst,
                 I => Y0h,
                 O => lzo,
                 OZB => FirstBit);
   ---------------- cycle 3----------------
   pfinal_s <= "011011";
   shiftval <= ('0' & lzo) - ('0' & pfinal_s); 
   shiftvalinL <= shiftval(4 downto 0);
   shiftvalinR <= shiftval(4 downto 0);
   doRR <= shiftval(log2wF); -- sign of the result
   small <= EeqZero_d3 and not(doRR);
   ---------------- cycle 3----------------
   -- The left shifter for the 'small' case
   small_lshift: LeftShifter_27_by_max_27_uid6  -- pipelineDepth=1 maxInDelay=1.2523e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => small_absZ0_normd_full,
                 S => shiftvalinL,
                 X => absZ0_d3);
   ----------------Synchro barrier, entering cycle 4----------------
   small_absZ0_normd <= small_absZ0_normd_full(26 downto 0); -- get rid of leading zeroes
   ----------------Synchro barrier, entering cycle 0----------------
   ---------------- The range reduction box ---------------
   A0 <= X(51 downto 41);
   ----------------Synchro barrier, entering cycle 1----------------
   -- First inv table
   itO: InvTable_0_11_12  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => A0_d1,
                 Y => InvA0);
   ----------------Synchro barrier, entering cycle 2----------------
   p0_mult: IntMultiplier_UsingDSP_12_54_0_unsigned_uid11  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => P0,
                 X => InvA0,
                 Y => Y0_d2);
   ----------------Synchro barrier, entering cycle 3----------------
   Z1 <= P0(54 downto 0);

   A1 <= Z1(54 downto 46);
   B1 <= Z1(45 downto 0);
   ZM1 <= Z1;
   p1_mult: IntMultiplier_UsingDSP_9_55_0_unsigned_uid32  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => P1,
                 X => A1,
                 Y => ZM1);

   ----------------Synchro barrier, entering cycle 4----------------
    -- delay at multiplier output is 0
   ---------------- cycle 3----------------
   Y1 <= "1" & (8 downto 0 => '0') & Z1;
   EiY1 <= Y1 & (0 downto 0 => '0')  when A1(8) = '1'
     else  "0" & Y1;
   addXIter1 <= "0" & B1 & (18 downto 0 => '0');
   addIter1_1: IntAdder_66_f400_uid53  -- pipelineDepth=0 maxInDelay=5.3e-11
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '0',
                 R => EiYPB1,
                 X => addXIter1,
                 Y => EiY1);

   ----------------Synchro barrier, entering cycle 4----------------
   Pp1 <= (0 downto 0 => '1') & not(P1 & (0 downto 0 => '0'));
   addIter2_1: IntAdder_66_f400_uid60  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '1',
                 R => Z2,
                 X => EiYPB1_d1,
                 Y => Pp1);

 -- the critical path at the adder output = 2.02365e-09

   A2 <= Z2(65 downto 55);
   B2 <= Z2(54 downto 0);
   ZM2 <= Z2(65 downto 17);
   p2_mult: IntMultiplier_UsingDSP_11_49_0_unsigned_uid67  -- pipelineDepth=1 maxInDelay=2.02365e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => P2,
                 X => A2,
                 Y => ZM2);

   ----------------Synchro barrier, entering cycle 5----------------
    -- delay at multiplier output is 0
   ---------------- cycle 4----------------
   Y2 <= "1" & (16 downto 0 => '0') & Z2;
   EiY2 <= (5 downto 0 => '0') & Y2(83 downto 34);
   addXIter2 <= "0" & B2;
   addIter1_2: IntAdder_56_f400_uid88  -- pipelineDepth=1 maxInDelay=2.02365e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '0',
                 R => EiYPB2,
                 X => addXIter2,
                 Y => EiY2);

   ----------------Synchro barrier, entering cycle 5----------------
   Pp2 <= (6 downto 0 => '1') & not(P2(59 downto 11));
   addIter2_2: IntAdder_56_f400_uid95  -- pipelineDepth=1 maxInDelay=1.277e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '1',
                 R => Z3,
                 X => EiYPB2,
                 Y => Pp2);

   ----------------Synchro barrier, entering cycle 6----------------
 -- the critical path at the adder output = 4.97e-10
   Zfinal <= Z3;
   --  Synchro between RR box and case almost 1
   squarerIn <= Zfinal(sfinal-1 downto sfinal-31) when doRR_d3='1'
                    else (small_absZ0_normd_d2 & (3 downto 0 => '0'));  
   squarer: IntSquarer_31_uid102  -- pipelineDepth=4 maxInDelay=1.31465e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => Z2o2_full,
                 X => squarerIn);
   ----------------Synchro barrier, entering cycle 10----------------
   Z2o2_full_dummy <= Z2o2_full;
   Z2o2_normal <= Z2o2_full_dummy (61  downto 34);
   addFinalLog1pY <= (pfinal downto 0  => '1') & not(Z2o2_normal);
   addFinalLog1p_normalAdder: IntAdder_56_f400_uid105  -- pipelineDepth=0 maxInDelay=1.20065e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '1',
                 R => Log1p_normal,
                 X => Zfinal_d4,
                 Y => addFinalLog1pY);

   -- Now the log tables, as late as possible
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   ----------------Synchro barrier, entering cycle 3----------------
   ----------------Synchro barrier, entering cycle 7----------------
   -- First log table
   ltO: LogTable_0_11_83  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => A0_d7,
                 Y => L0);
   ----------------Synchro barrier, entering cycle 8----------------
   S1 <= L0;
   ----------------Synchro barrier, entering cycle 7----------------
   lt1: LogTable_1_9_74  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => A1_d4,
                 Y => L1);
   ----------------Synchro barrier, entering cycle 8----------------
   sopX1 <= ((82 downto 74 => '0') & L1);
   adderS1: IntAdder_83_f400_uid128  -- pipelineDepth=0 maxInDelay=2.35e-10
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '0' ,
                 R => S2,
                 X => S1,
                 Y => sopX1);

   ----------------Synchro barrier, entering cycle 9----------------
   lt2: LogTable_2_11_66  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => A2_d5,
                 Y => L2);
   ----------------Synchro barrier, entering cycle 10----------------
   sopX2 <= ((82 downto 66 => '0') & L2);
   adderS2: IntAdder_83_f400_uid137  -- pipelineDepth=0 maxInDelay=2.35e-10
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '0' ,
                 R => S3,
                 X => S2_d2,
                 Y => sopX2);

   ----------------Synchro barrier, entering cycle 11----------------
   almostLog <= S3_d1;
   adderLogF_normalY <= ((targetprec-1 downto sfinal => '0') & Log1p_normal_d1);
   adderLogF_normal: IntAdder_83_f400_uid144  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => '0',
                 R => LogF_normal,
                 X => almostLog,
                 Y => adderLogF_normalY);
   ----------------Synchro barrier, entering cycle 10----------------
   Log2KCM: IntIntKCM_11_49946518145322874_unsigned  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => absELog2,
                 X => absE_d10);
   ----------------Synchro barrier, entering cycle 11----------------
   absELog2_pad <=   absELog2 & (targetprec-wF-g-1 downto 0 => '0');       
   LogF_normal_pad <= (wE-1  downto 0 => LogF_normal(targetprec-1))  & LogF_normal;
   lnaddX <= absELog2_pad;
   ----------------Synchro barrier, entering cycle 12----------------
   lnaddY <= LogF_normal_pad_d1 when sR_d12='0' else not(LogF_normal_pad_d1); 
   lnadder: IntAdder_94_f400_uid164  -- pipelineDepth=0 maxInDelay=5.3e-11
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => sR_d12,
                 R => Log_normal,
                 X => lnaddX_d1,
                 Y => lnaddY);

   final_norm: LZCShifter_94_to_83_counting_128_uid171  -- pipelineDepth=4 maxInDelay=2.17565e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => E_normal,
                 I => Log_normal,
                 O => Log_normal_normd);
   Z2o2_small_bs <= Z2o2_full_dummy_d2(61 downto 31);
   ao_rshift: RightShifter_31_by_max_30_uid174  -- pipelineDepth=1 maxInDelay=9.973e-10
      port map ( clk  => clk,
                 rst  => rst,
                 R => Z2o2_small_s,
                 S => shiftvalinR_d9,
                 X => Z2o2_small_bs);
   ---------------- cycle 13----------------
   -- output delay at shifter output is 1.71795e-09
     -- send the MSB to position pfinal
   Z2o2_small <=  (pfinal-1 downto 0  => '0') & Z2o2_small_s(60 downto 30);
   -- mantissa will be either Y0-z^2/2  or  -Y0+z^2/2,  depending on sR  
   Z_small <= small_absZ0_normd_d9 & (30 downto 0 => '0');
   Log_smallY <= Z2o2_small when sR_d13='1' else not(Z2o2_small);
   nsRCin <= not ( sR_d13 );
   log_small_adder: IntAdder_58_f400_uid177  -- pipelineDepth=1 maxInDelay=2.42825e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => nsRCin,
                 R => Log_small,
                 X => Z_small,
                 Y => Log_smallY);

   ----------------Synchro barrier, entering cycle 14----------------
 -- critical path here is 1.307e-09
   -- Possibly subtract 1 or 2 to the exponent, depending on the LZC of Log_small
   E0_sub <=   "11" when Log_small(wF+g+1) = '1'
          else "10" when Log_small(wF+g+1 downto wF+g) = "01"
          else "01" ;
   -- The smallest log will be log(1+2^{-wF}) \approx 2^{-wF}  = 2^-52
   -- The smallest representable number is 2^{1-2^(wE-1)} = 2^-1023
   -- No underflow possible
   ufl <= '0';
   ----------------Synchro barrier, entering cycle 15----------------
   E_small <=  ("0" & (wE-2 downto 2 => '1') & E0_sub_d1)  -  ((wE-1 downto 6 => '0') & lzo_d12) ;
   Log_small_normd <= Log_small_d1(wF+g+1 downto 2) when Log_small_d1(wF+g+1)='1'
           else Log_small_d1(wF+g downto 1)  when Log_small_d1(wF+g)='1'  -- remove the first zero
           else Log_small_d1(wF+g-1 downto 0)  ; -- remove two zeroes (extremely rare, 001000000 only)
   ----------------Synchro barrier, entering cycle 16----------------
   E0offset <= "10000001001"; -- E0 + wE 
   ER <= E_small_d1(10 downto 0) when small_d13='1'
      else E0offset - ((10 downto 7 => '0') & E_normal);
   ---------------- cycle 16----------------
   Log_g <=  Log_small_normd_d1(wF+g-2 downto 0) & "0" when small_d13='1'           -- remove implicit 1
      else Log_normal_normd(targetprec-2 downto targetprec-wF-g-1 );  -- remove implicit 1
   round <= Log_g(g-1) ; -- sticky is always 1 for a transcendental function 
   -- if round leads to a change of binade, the carry propagation magically updates both mantissa and exponent
   fraX <= (ER & Log_g(wF+g-1 downto g)) ; 
   fraY <= ((wE+wF-1 downto 1 => '0') & round); 
   finalRoundAdder: IntAdder_63_f400_uid184  -- pipelineDepth=0 maxInDelay=1.0503e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => '0',
                 R => EFR,
                 X => fraX,
                 Y => fraY);
   ----------------Synchro barrier, entering cycle 17----------------
   R(wE+wF+2 downto wE+wF) <= "110" when ((XExnSgn_d17(2) and (XExnSgn_d17(1) or XExnSgn_d17(0))) or (XExnSgn_d17(1) and XExnSgn_d17(0))) = '1' else
                              "101" when XExnSgn_d17(2 downto 1) = "00"  else
                              "100" when XExnSgn_d17(2 downto 1) = "10"  else
                              "00" & sR_d17 when (((Log_normal_normd_d1(targetprec-1)='0') and (small_d14='0')) or ( (Log_small_normd_d2 (wF+g-1)='0') and (small_d14='1'))) or (ufl_d3 = '1') else
                               "01" & sR_d17;
   R(wE+wF-1 downto 0) <=  EFR_d1;
end architecture;

