library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.Pack.ALL;

entity AIScore is
    Port ( CLK : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           Initial : in  InitialArray;
           Eta : in  STD_LOGIC;
           Result : out  STD_LOGIC);
end AIScore;

architecture Behavioral of AIScore is

begin


end Behavioral;

